module hbram_top #(
    parameter       MHZ            = 200,
    parameter       RAM_DBW        = 8,
    parameter       RAM_ABW        = 25,
    parameter [0:0] CR0_DPD        = 1'b1,
    parameter [2:0] CR0_ODS        = 3'b000,
    parameter [3:0] CR0_ILC        = 4'b0010,
    parameter [0:0] CR0_FLE        = 1'b1,
    parameter [0:0] CR0_HBE        = 1'b1,
    parameter [1:0] CR0_WBL        = 2'b11,
    parameter [0:0] CR1_MCT        = 1'b1,
    parameter [0:0] CR1_HSE        = 1'b1,
    parameter [2:0] CR1_PAR        = 3'b000,
    parameter       AXI_IF         = 1,
    parameter       AXI_DBW        = 32,
    parameter       AXI_SBW        = AXI_DBW/8,
    parameter       AXI_AWR_DEPTH  = 16,
    parameter       AXI_W_DEPTH    = 256,
    parameter       AXI_R_DEPTH    = 256,
    parameter       DDIN_MODE      = "",
    parameter       RDO_DELAY      = 4,
    parameter [4:0] CAL_CLK_CH     = 5'b00001,
    parameter       CAL_MODE       = 0,
    parameter       CAL_DQ_STEPS   = 8,
    parameter       CAL_RWDS_STEPS = 8,
    parameter       CAL_BYTES      = 'h100,
    parameter       TCSM           = 4000000,
    parameter       TVCS           = 150000000,
    parameter       TRH            = 200000,
    parameter       TRTR           = 40000,
    parameter       PLL_MANUAL     = 0
) (
    input  wire                 rst,
    input  wire                 ram_clk,
    input  wire                 ram_clk_cal,
    input  wire                 io_axi_clk,
    input  wire                 io_arw_valid,
    input  wire [31:0]          io_arw_payload_addr,
    input  wire [7:0]           io_arw_payload_id,
    input  wire [7:0]           io_arw_payload_len,
    input  wire [2:0]           io_arw_payload_size,
    input  wire [1:0]           io_arw_payload_burst,
    input  wire [1:0]           io_arw_payload_lock,
    input  wire                 io_arw_payload_write,
    output wire                 io_arw_ready,
    input  wire [7:0]           io_w_payload_id,
    input  wire                 io_w_valid,
    input  wire [AXI_DBW-1:0]   io_w_payload_data,
    input  wire [AXI_SBW-1:0]   io_w_payload_strb,
    input  wire                 io_w_payload_last,
    output wire                 io_w_ready,
    input  wire                 io_b_ready,
    output wire                 io_b_valid,
    output wire [7:0]           io_b_payload_id,
    input  wire                 io_r_ready,
    output wire                 io_r_valid,
    output wire [AXI_DBW-1:0]   io_r_payload_data,
    output wire [7:0]           io_r_payload_id,
    output wire [1:0]           io_r_payload_resp,
    output wire                 io_r_payload_last,
    input  wire                 native_ram_rdwr,
    input  wire                 native_ram_en,
    input  wire [10:0]          native_ram_burst_len,
    input  wire [31:0]          native_ram_address,
    input  wire [AXI_DBW-1:0]   native_wr_data,
    input  wire [AXI_SBW-1:0]   native_wr_datamask,
    input  wire                 native_wr_en,
    output wire                 native_wr_buf_ready,
    output wire [AXI_DBW-1:0]   native_rd_data,
    output wire                 native_rd_valid,
    output wire                 native_ctrl_idle,
    input  wire                 dyn_pll_phase_en,
    input  wire [2:0]           dyn_pll_phase_sel,
    output wire                 hbc_cal_SHIFT_ENA,
    output wire [2:0]           hbc_cal_SHIFT,
    output wire [4:0]           hbc_cal_SHIFT_SEL,
    output wire [15:0]          hbc_cal_debug_info,
    output wire                 hbc_rst_n,
    output wire                 hbc_cs_n,
    output wire                 hbc_ck_p_HI,
    output wire                 hbc_ck_p_LO,
    output wire                 hbc_ck_n_HI,
    output wire                 hbc_ck_n_LO,
    output wire [RAM_DBW/8-1:0] hbc_rwds_OUT_HI,
    output wire [RAM_DBW/8-1:0] hbc_rwds_OUT_LO,
    input  wire [RAM_DBW/8-1:0] hbc_rwds_IN_HI,
    input  wire [RAM_DBW/8-1:0] hbc_rwds_IN_LO,
    output wire [RAM_DBW/8-1:0] hbc_rwds_OE,
    output wire [RAM_DBW-1:0]   hbc_dq_OUT_HI,
    output wire [RAM_DBW-1:0]   hbc_dq_OUT_LO,
    input  wire [RAM_DBW-1:0]   hbc_dq_IN_HI,
    input  wire [RAM_DBW-1:0]   hbc_dq_IN_LO,
    output wire [RAM_DBW-1:0]   hbc_dq_OE,
    output wire                 hbc_cal_pass
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EsINo7+AIrgRtA2LbUaYH74B57yiINVyTSAxA14zAufIE0X3B8iwF8mscDHWfPFv
Ch/gOVeGjGAFtubZYvKuralSp84CBSTXRPMnx+bmWsmbwW2GNrUhGSczWFvV/1fA
ZvK3kjb88ZaJYesw9R66s/ect5lBI1nypeOB2eQvTq3urGZelDDloYns23zQyJB6
JyRU3ubO0LlcV5uECcxNTLxCl+nEc9FG9+q8a/qqYULB5pWSaIVFW4RLY9rfN69D
k9zPm6Uvl8Nq96ihjSDKEulnTrD1MgbZXf25NHtAG0vJBG2S806rvf/UJaCs0Udo
CTS+cgxbyYHJcJ6Z37jB/g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 152816 )
`pragma protect data_block
rBQRiZWApeIQ/TliSbtFXiXpYtKAjs3vKGs3d41Lw3/XroscKX2TdGOohTA84v5J
P1L10aW2J4S8IUAHG6ZWW1rjyeGz+dVWY/qhuEk3xbbPQz5MONG1X+WatOnKVXCM
Zgv3DoL/kvvzrKJpyp0Gutfl1tCAfYbGYIH5V5p38xvUgCg9GLzBrFFZYW++UkNi
jp9poqP5kDKKfu2ZJcQcXqGx94T7URjOr/dscfwTYrcUgvFgjK55A68mWlTu9aDL
0cpIAiSAPLCYGEr0UprR4v6jXv1HugWHYlZo+zJWq8GgqxnFtn4AcIUg4Z99rWCU
qIgQzemQlk6m9IVC36UoGLBwZ90cE4iK6a4MXqgN2m06Mn1QNFd7vU+hK/BSlNQk
hMkLyoE/1e3x0zmI15Jfz2wHIwm62uEAJOdzbAHrly9kaisRPJmBIw0l2KqxVvWN
R1NNmwn9yQzQBx3YIDAwue7KE0yY7RmflRVP4KRodY0SB9bsBJhz5xIkBRk3HZEr
gFhpg3UOTpijx1mkzjbAD2ljMlZxPKicMP6yQ5CKz91VGeGrE5zaPUiPc7C6DbcL
wOofyPAVvbQ7vMCuiU2o8pIkkn+lekun1brj+vG59EhFjYauh7lgaNkO+3tP0QV7
Qp1enrnweUA3rVy3gDw0tbhwxnZrvgIyfzhXXUgU1EkWNiKoOui17YIE8xRc7QEv
mGDGagj7O1epXpSQONOl9LZrknd/tKgSwr//kAAY1lsgGGHXMiZ3J12wefPvwoz8
sPHqTxJBLwooczAsQZ32zV0wdULnrUmRswGtEhxvdjn7Dhdb6KzeJOexOnmcx2vY
rxtLULzZMbsb33PcbeZewVqaAE0JF2SNLTJsaS9FAjrN76JOI4saRDXYXGCvxW2b
/+h7POuRXPEZW4chVJ1dsFbFRxLEMC+5MKWXLo9y/MNvmV5NaAzNDFMJB5bMxUCB
V7xAgREerjfXMTtG4+4298vRliqzOBGd6YCqLxSdenHcKRHBozCPjdOHhpUxjSUl
9RAvuFlx90uA5JSozZ+ny5fKfGEDCu28VKc+a1sDGOZxxfgYC8UtKoQ4ZcMu/ci/
/fwkaFugHfxvHEPEHO7tBmEBtL1QxniNfuhaWCFznjf5a0c2rylbnKpkt0IZv5SR
8Ip0izRmeEVhdjGi4957HVXkxcAXiVnbHjJLwdrYTsQOu+hH1wQuzZeftpWOPRGm
KIIokRKco9qJJxes951OveygsjpSNvxwX0sQUs2jMlyHHniN0y+RvbZA6okmxKLS
KMwI4se/YrydK0YgyPP8zmIF/JqtNERN8QLAVEKHg6E6/ID5yKA5n87dmt27cdZY
V0sXSMy+5xl5MxABHPGMvTtXFuJPJW3bmMVIUt5ifU0PthsBc+piTiiNJ+boMtu0
433zP10zMd7rUPljXgQ6n1Ua6uhVwqAC0s13J9sByV/aA3hDIDupbdYHUI/BFodz
KnwAjUfLPAJ4C08ZgO2QJg+cpODD0Ggk9UyOM5hwThDOlVU5wMQJbdm5UVZdFBlg
7BPEZCcLPSjea+ddKBTfNQqkaTIkJAlRhs3zj0/9BZKM16+tuQFCbFpeL6D/38Wd
LUfqP3tIAqrE7MnNGrsMxD29lb3QuGDimRQUVanZCOB2NmzYTut+EtEbK8IalSeu
GMPGZmjR7ZQMtfejAzV9ehPe+UQT90U9WPReyTopdVS3H2gB3SCxWuX6kDsZDOvt
oxEL1xjck/uOu8RTb0BzwPts86iYA8M2JnS+24Y3gKUoZ0J9JLp+1k8Qj7nmVGtr
tCNa8a7J4dNbIBAeiURexPhldhbEARXG8egS2wIXB8IRoseEeFJtBcL+544XAu7r
vEfzKkrTABskFs12EKor9YOCSoYiM19PazSg8cjcNqZLf8YG7CHbB1ydbvGlma/c
OKH43xuQxVjbUVREP/CAzMXSbSTpuAAkmHMLBrDY5GNyKf+sOS3Bz5ixsnYUFuTw
CSgb1DuFPpCcd1+YZ6Mwsd0WfIXk6U95IJ1YNHhL8URyzFi6IXg0f3PAvQJ5m82x
ZkcDjZBv1M1v16kj1Lg9ZSRUZVojhhkDETuEzmVyt4wqjMYdbnq0g9m+fJh5kCxg
U0yhHVT60SqL+jQSwDjv+HfNhC7l8WuFMIH7dxu4gGVYWRGkwHuDrJfIe6KX2KOl
Lt3ob5uczdXZcPzkowkb1F8r/T7OXiuy7fF4Kad3NaioDpVSezJQkcgakeazt9N2
9J2sTyz0jzX7K/HMj+CMFKUu5twUaODQU8vOIrhG+tljgC+3gbr7YtA5SuAqSktd
otlxtIGtNiADeYzYYPEPoY56iYr4yLMoQ6KXMmbp5DYtBEk8zdf1FefP7JL/ypky
ABRl2NPDN/wJqfy0S6f3kRyqAljF0SWt6WipFEE4VqPCIt8KwlEdbJ1xvx8aUWgc
3S2DLR+/xjith2oiPr7FrxrRYnXtqd9WWwmdA9h+tvEiUeTgrWuigCCn8w/cvBjX
tfO0J1PFQWCHzVhv5oHjFCKEw5UccEDGU1aBazE8+s9rEqfoxMZogLTXhQVKWxxu
UNpP7rSVIyMhbgF7jg15zX12wlwGSfX1HFLsuPU4Ww/EQ6aj7VZyBWnXTMgH0boU
8vef8QTaCFFIv3ax6pt6IV9S9kEFdCeU89Ea5wF6MC99ivXwflqXmOS+W1aTcQhH
oDIUminOmvXaHmapMMKym5iIF0OSiJXFJRHVL5jKsnBC/4P2X8pSiG7EIy5I4FTP
ApZNi5TvJji2UlAKcQBAOyJJcXGNxs+UL4Mz7BX4JV7plQ2tCCBjdoF4wPs+h1Ql
Zdkr121puHxi/WeEscq+nt18m5A7/VMrqZjOmw9omG2KvZnoiqcvECVXiOE4/GwP
IeSntblSaUo4oO7LShTTJy9MahrvFVGogCuGp98gU7PD0weT3KyRorrsvfuZbDxS
8w6mpnzfj0HEnDaAOlJ5K0DkkAQyzPDBefjnWfR+Ib3/jOPa2ntmTqd2NlmnxKoK
uKMJB0SSbjKMFGgoyGaZUy2HR7UMjv8yDJdf/UA2801c5BJhBqakUUm/FsCdclJL
Ue+En3ymGtpZcVG+tOnGWKzB1LlLJz+6LelFaNXDaCd2qXZZXwJX1nDwMvfCBJRg
Pr1XaKHwlpfWqK/Ih/uV8sbJZzfibXFiEEdiOaRaui0KNew0TI99F3coUvKJQAyo
Y8vZ75SDnxqE3LW2Wi82+SfL6WZgvsu8Qz6uISw+y7Z/HByvd7BRUkrika86Jo4R
c1tPcBSZ0UuSbREGqUzugwyuWJiU7D3DYyAsACEH4bA6xkth0W7439k7u8vzRqBt
xICAtaBhkAD9VTxT1amteoQXSukdYbaANI5WNjcVcolg3BlGHtAcyB1YAkU23TII
PkCEnkN5BFGDBvakjj73DRTZRDuDMxnywA4Aih9L5CradYKE1dqklqs27DMCvGnc
4zV5u6n0LoRVGrYGqYeByCzTucKfTAwVFQrALC29ERt6L+gbRvenC9ZT0MXNhxLi
Icd7jcfUNOZOK1rhScn3CQapyPpr8PGDWOSYDadnVo4XFo5oJGRMNn4W6PhHaEps
NQi/ZkHOFKBTQlSWQF/YG2o1OYn36YszPC9p5XqW0SRV/6B7a0PC5+KPACbqB1bx
/Vu4hnl9C13JfJqsuOTCWlmPTok7VZv+cEAnh1hgbyKUA+ybQng4XEPOIgyHTeVJ
KJdSLZ2vXo3OU/BHflg7bhEM9pjZKP+mWztRlbaBCaUgyQNQ+P7wY6iiofsp6zzy
L1aUG41PXBFJSlixiBukLBtrlHjeJAj0ivZo9umYEWR0bi+4blxtmX6XfUNDVP00
RplpFyI3hE/PDcP/5HqL4J76BqzP6KcSjEkUCDwZVLpmLLmD6eHG55f7R7d1POpm
pKhiLkVV8VYzKzzwBTQggOGvz8PKnv4m73pr23AAQoAKgKhp+qKPtn3EYbKbp8NA
AYrC7Nps4PH4MNftvwgzGv35LNzk0OJ7s10Y11yyRXuj8LxQbbx46Gzza7dwnobO
rPa6J7ximqY6sQKBlg0LZknW9Z5/O6DX+1ilatTcs14FgruTXoSkQQlgqza7GemA
MIOf2TTQbMZcvgTo7gTvNMtf9UxPK3UYSRsR1wctQsl3CMxUSKgC/07kcI3hn+t5
ScYZCSHLRFdx3cAesLr7CT833ZEAaeCoFlcxjCSctEoTPqcPbOVmfQCVMe/EV9RI
In+8Y3WQae9EtNXsYikL8+e28++3bGu5nWIHS5cq3YTf8d3Ht95xeso/llaLeWvF
bCRiXW8QImBD08Xl5andIhmW4yLP/SUpMlOujBdpwQHtbRaPlOAWtAy7FAlujaM0
0BNXaBiCjPjPvmpE5mKaYNqFKUIiO9S+F8uQO5GbOyMB8mxckGDZ7G74Ye+rxwnB
hKWBqcsOS+P0hUOVXMjJxJ7/gVNVv4VMZatm+XwG1xA9kezODfB+mPhcrchVsy6V
wsDrMqayAkj0zauBLPU0tu1vJfWsBV1bMuot/JKerCOKttPYcuZhBcJVFYUF+04U
7WYS+8yvF1JszlFXRmWdCXTtYAhQKNvU/hV1Lfouvgszv1fQQlTgJoXNo05DLyWa
fXV9ZEb6AcCH2nrcJLnTz2AxTrhFfth+Mh8MLfzxbx66oAfbTy/oPv0G/+GO9Fes
yD9QHl1qG2P5HVB/6eN8eqQLjm/elB3pEVEhjgpPo+8e47cwi/igwkpzoYF9dElW
9lXskMUJ0zcATs4mpM7wHNoaD1JwTl4itHFJ+KEgGUwlb+/yI/kE/A0MtLfXmAr3
iSKZpWPuSo4JGnViaA8X/1eoDZz9B0VdywQM3wobBSxkoOwqY8f/l+amEz5Fcnry
n0gWqW9VnGhTYbIWCNoF9+kfsk5hjAsRBTU42SptQhmuXLrZh6FIfoatopQsYLuy
8SQKaYt/G8+k00Tv5Ox796moDTGr9m0iXVY5FzIcLhegv/OuVEWFvRuHB4/kWXjM
xGH+xnJObO1LD7m8UyArdVk2eeMAQ0bKV91CxCqU/wTtqHVJN65Af+Blwnv9ampr
pLVzGVKgrGh+/Ijkmyr5PT0T6yIP2VrlAMixrxxHARyZLM0yPLgAzNNJm6PkNqM/
jzlG5Qd2WWGaOXzyhMCCowX0rgVA1XFNYhRZHAB3LrBveqQc8aZjYL4yL6zCsWlV
aecXvXaaIKfNc2HQGuecpPlqK/vR6S6f7remi+7vgCnd4xZnVLd5bz03DAtXTw7l
y8uOhagJZ95V9xeu1kOVdwZNjwJ8wmRhA0fOLaUwrb5545MKcjTszhSksZ776iY4
YZYPXLf7Hen99zKIGfhIHTzm0HQ/4v+8a8c8KdV8ltB7asrorvj8GsghxPiufe56
JTWeQ19FSYwoEPQaNpxOlLV4V1DsBiuVyQyoRg4IogUl7qzS+nHDe0x99YnWQqne
x798/baMRoikYBQ3pyv13s9gMdeIWZ/NPLocDW7tKYqvCCvhtK8rE9YAU3P6Iel2
uF4nrw4aowNGkUfE9zIkb76fckECq6Kkh4Gj7pOFL9HAPAp7jZiqz3xXy8BqoLBj
0pZUR8i8b3B3j+tJicWL0fq1avfD/vnzXrMgBo7yUC1VDVlnzJxossB2BpChLwo8
cgUG9aN+vqO+1pGqBYQWu8CsfM1mEuW7qJu1PnP8JdyNEBO3a+QfydP6TBCAS0CD
qhneb8DS1pUlY1pcs4zESPGHtaZrmdqIcZzY5TBkIpXZOriZvA9KjAnI0v+uEp1O
5BMrsgx17ZqaHOOPOt9iKK6mAhaerxrBo7Hj49A2rxvL4q+tPFQYSMRY57AvoNvt
CDEdzza79UH6byIQeMnds1nJNH9o8YOhFcpLvpUC6KHdgrmjTG1ST8spn5C2NXo1
mdMGz/GHFrdXu5ia6Jt5arNlgTwToF9cmEHIm2uCDpdOFXHkAlOOfwMfNhTFFnvi
JiwKVCCYE1av6X5VTKL3oZmTv9xtpL9iEseMdOofDrXKDLnRxu5b3ekx6NWVF1bb
vV1SYolqpkR2nud+l6/JKDw6OV4FnwcDIB5P5BnXtEyFQCgx1TexiUGmwVUTerY6
Y+XUW+Ipoh2sBIeElrmRPztE8iX2afPHTcIpz7OXzzmM30UBdYgO+IwqhqFx3kZh
wloJkTfvkFhi0ztC62WKphClZ+BXEOdN1HR7O9vhJuxsp+8d9D8yfUg0KOhHa4Tk
Rey6hRWOms/bbl0WK6i3VbNi3LzsND0iydvrIa7pY2GPFZIFj+dYXXXMFaNqjR7D
W4rKFiwliH1mcU8P79gVTdnVB7vYxtaRIR6Zbg52mbIN925tXZHFiIXWjvOrjp0l
qasKNbDNOR98VMa0XWYPkSdFAH3rfxl7fgsI3GlYYp6wj9bQ8M47xsUgzuDg021f
1nuvgnzMqP88c7faf60lQ7Ei8CZVk+VOYblLoxRXbGyJsFFEGOZmUxQNjfPfR8lX
Gh7wJxgtbCFlCCes9U6s6HqzxdyVlCmJQeAU/Yc3lum88EjqjncfQBiNPSSkkmv7
yNKoN/Gb+2tVY5nSYQiCG5WLn5bDWt2THcXn2G+2MAZgWQxRVAxfQJk0V/RAPBh8
axgeO2xycmLFyxACSlFQiefS4W4MpQWOXBEPbxViutIBa1vhUskkwRY0KvvBDTxi
ccaf2Kt+qKkKqKEXSGqQlD4gPWdDea8glzwHzHP8ylmg/2/tPfTbc5NnLckUbzxR
pjWTbQftZELq5kpLWoB9tOozjKu/YEJwzyL+EMEmMSJJkwZ9s2gmookLD+aCkCdZ
YXBdiLPUxh2HOfW9vnuqAgGvjzSyvC1KJpLHOrlBl6CETAk59XQipsEL28EK2n5x
aZuUR8u5MbiaDe7PxUcHxAd0Gb2BpaJrI8YrZrMU8Ffto9yQFktl4xKEBiPdiZr7
1tKCNTdIov83R/UkwZS0IpOFuwmzBpf0IbJNQMxMBXoJSFPBPQROirvLbunjQXI1
ROPFG1Bf4PriUaO+OzVtnfNTkEUzL9mLl0RPvLXBesoVYKgPi17zHjEdMHCR61bM
K5DVEblQetYt9umHcfqwUEEO8TmPzNcWcPHdjyWoVKME6wqvIqaGRc8iecXZF1CY
P3bZ8nZ2ha3FsX+hvwgyuG1HbRXkWO21mlzJiJrq/AI3+uNDSa4xDNtf4dMRywTl
ejcXn6Z2WzoJYpyj2+CJXNdnZxFCERliJZK9/+GMrLURnp4hSSJ4kNkaDBo6qXdZ
5RarccFlVVimY6G7e+Gv2MDennEJM54mVPapUH0yKHpRJOT47pqdHob5wZADWGbX
Eq2hnzO8T5byHoDj2SXM873VjW201KqU8o4W4LojaQC2dVwo6LUkP3ke3eE0k89V
fTu3TbQ218zth3iTghHoWGbGav1ZVJ9fEPqnOtud8s3Lk2u/Ylqofiouy+TcF735
PFVNcnjVqg2VBUpFSNMI4wIqVZ+EO6v/FkJcwAofOxcEEP8epWzRdjsrZffAODuY
Z97fAp7DRm62Mq1efuiAZOMEkNf+0S5FLxFKmAxDoBoR/a/qMAIE2RV5oHpcSxhJ
3BAcv33z02OL8B0FBgyWQK1hPZxV1gjA1hHwQtmM1/QYw7pgAZBsJh4mqr06AUJL
ln/sc+KJXFj/BjG1iyC+8iW+uO+VWrRjK/EfrTNl5RsyHI3D/0AwJdlT0NmOEjgl
YAaotHOGfpWeI6fGLkNhZ9fEHgJuwV9BWKLC/3TKGYat9C5T9Jlf7s33TITOYwxZ
xt2GnLCu7p5BHQHPFyJ7UgwYJX7YuIQ7hGLPD/dgMNH5Gwvw2LC19DioxTpGYSgA
LZZ/MCoUHAG8VFetvOUWfhkqIPnJ5/NI1OH1/qleH9kjLPm2rLFY+G1502sGFCoi
i4zrJK+Wi/luXwx4/6z1V3718klj4FdPbDcEfLS7HnL2uaKVBtYi2AR/HS1NC8mZ
E4g6qe92w5oitR6uvNPthNBprk8eWoHX2ZqiIdcAGVISOP4y2aVsdksgj/PaaCZv
59ROroAn4JQPlBia3lWV6YZC96ozrnbSFbValfM13Q/g71Q9P8GjkSRysnk10Ums
lJMh6ABnv/0rYISbW4bDz/bfQN6mVAdGV3Tza77K+ckXxrdu0Jd4wPLKPvufSnKD
KRf8Kb7e/kW5RMpakFuP5LdFq4+D2AhCvRLZUanfM6qSTMAfrR6rER5D4bvlXW9y
mMyPiJy/6HcnqmOdj/19/3EtGJay37ufebYt2nmwQVPAyHRtdVbOmGkU14cFm+6T
X9M16Yt52Kmtu9QKjw1J5JdFwOI45h1EpsKgukM90pGa4RPik0dUog8XqF7X4Jeo
AHGyWwjlUxbF67RX//jWyFmv6mefsvpdViV39ij4ZAppyaQU9i5k6pygYyAOBGNc
j7VgZfCAMTU8ZAokAGkc5NBFio4ZY/JkzJYIkcqXYt1xvixCOok74gcrBlevngvr
geeta9Byhc0a6B3hGdRqsuzmYIyPHnpH/eP3MqMNGdnL1qN6SUkQ6XkzO/b8hnz/
WRbWscNJKP/AZ6lShpdFZfvV6lDUXuZlIHBUc0ggx6IJTTV4827597IUJ6iYDVlQ
Ub4L/DW9myYaEXVbusNvy3PCz6p41oXrFEmLo379APvXBA6H7Qi2mev2/ezlHUrz
cBRbAN4Xm22Tqa7HIIvYSrNIxK3zyacAA6nfk63uUOtmhGpZM5DAmB01rnppZw90
33j7dTtueLZejx+nI6cffaOZSorVJ080in+SLyk+w0KwXYnl+BygRXsk6BkZ0Jut
J3nDj6yWjXcXdLYZiaJw6lKPfd+m5g3b3Ptonda2gGd7T08Qi8o5M8LYRiYZQPe+
TRXIH/eFqUb0w2nDQGy/ipBtWUpfJMrsqXOa2uanVHTeKVZvhLQKAA8d+YQTTDPt
T6RGjHkKkjzLst6L1TFg+G2jELU0nPqiLGDag93kDn92Gs/e9IOcxJPVZ7wu7OfG
hfJLIrX8eEoN9alhBzd2TOGrHJ1eo0SLLyfa3+DUNPlcoFqEqt9zazWgA8Netiak
AYXt35RZL6RBjSS8Mh1O1u07S8p6jVOS1T/uD1f7n2LGOD5j7vyuwXtvz7vfHeRu
xiqMwf7XlM+6ZMNkFfk/jImJg8Bi3e4nVvvLqEVbEL4HZc3BE0drYzuB8p1jhn+X
9FS2cL7UHzKCAJAoeR9v0l6Ryc0yCS1vdODwO/ZJ20Ss9j99SIycMWX6umSKkE8o
zzWGf6/3Zvn9Hd9A5e2M0VT3nSiWZpsC3DtP16LbgHzjRFkBuTAR/x/MkDIGZ+bF
nwF9fYqOjEl7T5hK1CM5x3FlmoA3QV5Av365LO7o2o6SuPK7hex3QJc+j26ENRkf
71CIIgYuz3JWHGmWfTn3fQpATMxdFIA/gx/bhyEnMKF7+ncMHVXHHeSit8hyWktF
JW916NQe9lV4ve1oIskBQV0f7HJh7coGVtOL4RR3LCItC+IxJoA2vCck8KXmGui+
hsDCeho1pb8rYYyNdFkO3Q7rzdZ70Fq9hHCbizB1+9aH+KE/SPgwNd4cZPyiugZf
7/Oi1WtrlxCBGynr0IBvC3mZGDmWfuqL2XGO93yh9HSmf3MF4k19Z3VnRL3N77cf
yFvQUy9HPbklJ3AzmbFRqvFvqZGC1L+amXaSqidSzpyrgjEShBW6svK1PJxJz+ev
WK8oysfEuatMSD4ymQOHgf7y5ov5I8N+6Yh/XwkDySweot7+ZmwNVfkCRxgUW60E
HewmzuZMcUtaxm/OmXsRnyyjjmGuv+n0st3sJJOlqZeXmblPZm46VyZang4nuD5w
VN3YWIm62AV2/KBXoVgXoi74Y4Rm+8UEN1o65cqQOLoV02t1JeaMrX2HbmamZa/0
QLoM4R8n4i8XKo1hL5EXuMtxNh/8Kn2vGJr15mUyh+8pcZjJSuZQ826n4uyU3KM9
tCl6UyyOatp5yezfWU4OkU51zI6N2V1SbixT9WV2Vp8y1K7WP6YNWnNzDpy+Cj6t
1+4iMncHyZnuohNrtfiZKjjrebPaXVJgLFqZYNBv7lDg2gLtCx1vNt+FQU2YvtwZ
cxAED7R5OJCial/PXFvoElVuks5FwPC6DMYmzLJ6FX5KbpCymV1/eOBCpnNyiDat
1kxTshq+NH9YOnQ3mlFIgJLWeUn8W6TuO6k92YTWkdvm9UoxtF/eIqyf6iScVJGt
FHMGm9i+zVYdY9bb89NDIa9bqJHhlMxz6I4lzTPiWF/mZtAWFMb+9gtDc2QMdKnE
jOLdojqbBIy+D2wq/wThgqZnbX94Uf4AMsNSoiAoOtTjOVQ7a+tebPWUqpVcfROm
vwU6+2ckbdXWy1JLmquBUl6MsGH4ia3/760bmAVNG8qUrQma4MxC6YDdsEqWcgiM
XR1qL6FD+JiowfIaqhaRmzPePQ3G3oqxklR7meW9SvRctELzMB2WX3J6319/qncv
iG2Gt+0StjNGCHG47/N7+uzaZ0DEO8N/ytU/Yz7aUheHehg3nSdWsde3TZtCzAYo
K8OEYANsGM08b6I4xZZs79RPa6UssSM2jdsR0m8tYK+OqeoAOppqqMKD/m19O5+G
UzjfWbamTexXlo59B9lcE0nHYvX51SV+LIBIo2OgYHGlQOEBfYJErWShTLz+qpVb
vu/ZfwXMGsRF6OYFOEKVZq/ETMhHrnad/QoJd4RuwASLGUvqZGosr0NWh9ySVd5p
3d8Ml0o5zdwK67gHLKcdJAeh69mpGeZOlVveJfj8Tqbro85LpIDXkPpDam1rUJY7
0VAorr5hr8nvvA9u75BnqKFi2c6sFF136PdaVCfGQeuGjSZ49KedNeZLR7vcFuqn
TjGYb43eVjOzR5fqJ82fysweGGHIsmjT9SFGAgQjKveWrDiqF9RpppAoiX6mhVkq
9MibRdUnMlJssRQuixA1arww9FjH/2tkoU3jycFLwJsUKnC3kV2A3FxIspv+Aypy
L7pl68cSuFUpX6lkSt+yMYXYDXicsHgt759cZa85ag20FqX02Y/hEspEALCVJ5DD
RSd+kaqMST0ItsbsJxhL/3j9LCq1l+2FxOlk8xQ35HPAKjYl5PNvnuz2bnnmmabO
ENuuyXUDhiVFqKuCvsBu9AH3sRc8vewTWQ9ANhPfDL3OuWYfwXh8IS+uCeLBuV2U
mtN+peQDWdm5WMvPzGchg3HjA/Bk/X/xrTlwn8Cns0Lzxhm5S0hsbziLsGY2Bf5c
hiN+EE/UbpxvJjZCL6ZdIllsLAPoQJ3KF9CPSIR/dtGR0e7dRp+g/6PPAcFcAX2T
n4dAIrLkx+7okKEN71KjEU+Io8zED0xcL9I7YeyK79ofBU8XtJNyWVrumdB1S+m8
1U5gqGp6+MVs2X8iBNnS4Xj7qvMj9UZqqQI79hL4BXwSZEgMmZh8YlXmLu6Jwom9
fvpupIOcGEWQSAqVCdGQJl8itoTJVjVX+BZSdAVOdcsXTX8Ugq+6/iTIptFxuH8g
MftgW8Evn+bSGr71eoJct1uJcutBDiKsFLR/aPduaEMDjD2jvLMUyaxPv2I24IG+
RnkgQUZCgTRaULVKe+tAa7PVOv0gIGKkcTd6prNM75RIDUevmAh7OWwmccp7rwgi
JB0JBA3uu3dqY84q29HoBj8UEV9xE/ugBr+3Rylx9zW4A6xghckDxnDHCcmr2esL
ufS06WorgGWVOkLbDLMqVZW7ss4pheYCIBoBWw5pccXnmSPk2oKQrrf0BsKQSOEu
tvsDqJ6PUWUTqpp612/SkMzCEmSNxy4XO6ve0mVdk3ESRJZNhWaMMaWoPbgNIIGX
86iBWoHBO0WJsjBPQ/cTWBIu+6VvoBt9CnOihaqOg7oZAA2+Vh7XHomtICc8MujX
59Z57V45LEtqE9pzkm46UGcLvTt9KYTmrN3dRrTIY9Is7zIWI3Kkpf2DIHiLzYI4
CmLORpLiumS7XmzoNIBWsGT+UQkWfpi4iNVPkVnr9da6l6Ow2cuyYkqvMYabjRCF
Sudipxqx18w3ziKkc5NzsCSzT/H4i8YeOpkQCo9wGwKmZDvMZyZnBSA90VMDxVmZ
5USexS77/YUISjEp7tuAO2TLwl8bRSXtpBDizF7aXjsV7HnoUeyxvQbofSFF6mxX
MxQv0fgvU7SMgGY5LhK5Zml8vDWzBy0yZz4+wr0KOezyfBulcHLLRMDKQDAsf7yL
d913lpcOw42Mdn4VEIcl8Ua6V3C0hfjibJ85FVeoyDGciznj+lMhOpqVB7oKxCde
TnXP6UFb+PX2D5igNv/GW3svFJiqoZ85Uqb9Y7z2GNeAeTCr9Q1GkccPcA0Rh3fZ
TP3XC4ShoS6AWve0jJ14yVovlc6NwhM97vJwEYoiXX1tJzPL9XfDjf0tk3+lQRAF
/kOBJi0+XR+97NAJaK97ztsWfTwPYTVdmX6iCZAPHlMiLq62xIqRo6JSEXFDsSIE
AeGZkLvrD4xViQKXRVV4BNaeyyD4OSDL+Pytp5b7lUUhIGMaFZeJrGZqAS3joA/a
/ThimKZCh9MneRYAjN5BTtmJsJirShyXdtNcokJXce5vdEGlWyv6Toskx/RQeEVH
syas05HixGlxoq4hLKD/HqyXqaRFLKPFrPQvZmknM34nl8aVGtwuj1VcI4c3vclH
YPP4eO5dncNN0I8LqFQFlSGDocYlj64y1J1NsUTcLq2C/yueMSnen2IJU+TMiZXT
qBrCHrxxrcs4zLkDbHOaKlcA3tQkVWD+YZiQ0MtYJbvngL9mcNPO/SgGA298fiLF
ob44TV76bm5xs+k2wPQxi5ym4jtp4JCL/BRZookyMlx6nuDz/P3V1v7SSx3nnvdp
0bcpFK2ii2+Y/SDl8Eh/9Er0FhoRdkpToc4k1g8ppJJkW6rSJN3+uugZH5+icBur
XclOnxFW/jvtUFU3yhHnKZe5l2nf2FUiWbz+5mrk95P0mCcQe2B/Tkr7Mg9g7Qg4
QvCOTeEXlp31pt65ixfhH+VxKZAivhuw59vJCQi0SWuZc5p6jumYPTnOuAXv5hCF
8m6xolbj3izbKVbcuAIsP2uGWquKmG7kKcMR7Y9Sp5x9BtIUASKvnypCpMpONesS
FnWr8mXjik/djocKEhusi7RCWl4+419quJ5ANPDbV6gYgq8PmoFtknCoD1HZoh7P
l0fceIRtquVgZwLqO1F15t2IzoGheFLtFkmWSJkH1aDpVO4j0zT+mDsM49mzKToM
xbUskYPiH7aYKdxHMtndeTKy02KPJ4xP6yAG9eHaUYIX6Z2eJnNYkdJyRxnpE5bC
gSt5DZBK7mRMS+bg1k5ZSJkQBg7HD1dniDG+YOLaTC+433PePRFwI4M0oUoPIZES
7ofyyE3bMIqZ2fC3MNG52IioqAplq2CfyTyY9WO/gi0E/68MCv8pU5mFKzook+OS
jHI0WpijaTbAwmTw7FVe/mlPhQVCZr/+x2IrGcTTBamTmeTKHMGiRKXFih5aVRmI
zsMqj2TLbG/rCHnKBmXeN8JLaSdYLUvdkM/GWX4ErZD+pKAAKwV3SffkkkE/vHvF
0Wx789ahnDZK29Z5iRKRnDpO0fJj6JFAbJacYrpklyeTSfoiScB15TP2ktyv9Nx5
rFA9902yErXkZ3s3tjqmIH6gVy2JPa+HPgOhvO0veoW4JXkNzgUdwV/8l5bDY8kx
oysZbOkFDYVbuI1i8ATjJkM4HkflYQLB/+sZdE21YkIg9q2FiaR3FOOGSzug4R6m
LczC1M3xXnDlCymLGlaOozo2RTulew2VaJJBXKsg0I5NeIRycLJnLiDaufFEYs1K
LfuDw42VYT+ZxxtmHJ2GjraEg9WNdFeocMV9660NPF/UjRvT9Uz/mRWAiT9Ycl2L
vyp2EObmHlb2P+WXrkX27LmkKEJOuKMOrRfgOoUNx36B7DL6JqUCecxAG/UPij70
9YOeSfPEjqSMjIeroVtzljp4rO9LFIs/9kCGcrc03HEv/L3pcf2MNP+Htt1vGMSZ
u8tDDKiakO53IvBen0Oq6MkSdzdUcY1x/z7Uq4jun7B+H9mI92q6qBlHG7blnOtV
9KAF6tMS6S2Un2wfex1DlEg66qXutMqK6Lu/imqxVseUjdtAJ9kRKFSgF6LxDdrg
Mk9B2qMLQpz8JQHqx1lZXTeWFvAXrLua9pgpwhFQaWSQ8lR0rXg+6Zxo6UQydLku
bCeMNCJu2NKW/tBxfVVxtH3csNV6e519Q6MNIVn8QRBF2VXCTEkW98EItPLNWd+z
o3QYADTkVsVseTK2v/53MRW9kPzLHGDbQEWLBJspanPJnOc3Qgvcb2eDUCKKqcPs
zut7rg0JxvptCgi1ipsE490hEWlOZjBPxNZ+7nYkg+d4HfFzxIyqdlDeqIMaH9TI
oVI4T0poB9THubtXgVizosAb3t6qxvxjrQSqxaX058EgPdm+utIqa9XEppOakoWS
MxJal9csg+JwHnrD5X/6absLmFQK5b+SiT0aE8vVC2tDaq32UIzgwXFnIlaD80tH
FC7i4hLOXDX27DlUopnRpE96LuxgYCM4EyjwOd6+IudFFjDtBmVDK3FMf4acH9Ov
BWRdd5UWhe2nLbQht7hFxkJbRojZaHGHO7dekOQqXf0F0DIq1y7fvYIRX9ODr9jw
p+5dCnDNJ9lSb7yLOTk2Uj7n8qTUz5kAs6VR0RYaURs0+SrgJ6buJbvkqO6vnIcZ
8u8eDuf7gbEOwT31q4YXqbigIVQySV+iq0QkIzjgWRoOOeJo0Drp0g3Sf4/Xa80k
+pcG6ox5UmEZ6gTdXXT4yJ0geVxi6n5ijZ2GoVRnzG1xO7/eFAeCB2Aj7igaPMFk
/ipDuu3JXKbEOEcdQo+XAsXjxSICJnMq6onE/jOx79N8MUBoagX5N9Fnxj4xt8s/
2iKem1yvZwU98V1lYo0eIUDlhRI0UfgL2OMFeIl9qRVh7/K4YAqpLOyTtijmtshk
UcQxyZsC4S6kh4PpuBa8OLO5toyIl14ZnYNr/hZZ6Q7i7Fqyy2Wci16StzmToNbC
60RTaIdLdOdb0ft9FJ1TNKEBzFO4n9ef+3NXcyrbp20rG080dpXSrHy6VOS4pdSJ
W7+F0DiSjxRrsyLsUQahDTdcJ511BBixIpKbZLcFf1TWbrHnXOAgauDlmiQH1jHa
BcjpUeFlrcI0KRds+mmgWPjJppeg9nbOLUt4KX8CpzmekvJ7UYWeQPwRbQugQBnH
441FuVPqrMpfYKJQzvN9JR8viRarfzP++iLFkBfk18L13o9SWCtCUpKtE0YHFuFm
gJBGerId3KUadWa78dXJYxCL+oUHNLKlodkmpgOVG/SVI3Oyj2HCcY66S/1Mb0FN
zoEZ5FuqH3asaAOK8MQBw/6wdr0SYcVUlMuohuOYFMzS+yWgAbsL98nWYSmiMtzh
Bl7AhhFK4J8xk8F9Xg68vihbd68WdFelEhC46z+EE4yVkvavmqJ7+oyzo7hN5dkw
Z9vRwUIRkxE8yps72Ddw0U2L8yHobn/aCAHR4Q16DoncnHFwCnWiJDfb6wQpcrHt
jjFTUImm1kJS/JrPKc9sKFT5hdjVuihyzLX/bagEmcsIST6M/c7Fhu0Ggv4vYDWF
5TRGjdfk+2f1n3IEUlvPMEGbvrxetZX+b9pOV5KfL1az4mwh7C168+5H7s96xqvn
3UpXNmar6mdxZKvkrRUdzpE+iw+UZwxrKzcsrwJnaiD79jlJAU9s4ojbj+HwBCkL
KE9UlTqA42Xyy19NoX5AHecwklKJGyrhha71yScgWq4zc2rTZVGk541QI78yrsC9
FKLJqfTYggKMj95luNUsFb9nccAC0bSR89Onx9puk5nO2KmYbhzmKUbYmi5vvUxx
LlPtOS4yDR+WcLAX+q+L4wy+jNCJekC0EKT+GajFazK7A/uAhcHlhDoMJbs0y/fU
d+3StNYJujSEVqSQvzW1I/I6oH12GK7Nf7e+eSTmtQc2eom6NcJd9yKLvPaWeXgr
1bKXE1C3csgSTYAM298Ce0iRCRc/+fYZjCIrb2D6v0lNmifyLlGpPGqdur+TFOjT
lvNVUgoexKikLjP8NmdHqBEVc1wQGkseK/Et4EAMeWh4hSWvLASpgpXLcL6Wlv7F
yCkI7OaxvUG5LsrWTBrt9EparJVtbLV3tkyOIkE1sH5VCMejLP6h8wxulznwXUyV
0Mij6P8vIFZCWKwNkUmfKDAkY8lWu188EYfp7fhFZCnVgejlyUlV/tjWS8uXvYQB
aL79xY/cl0sn5uIUYBh+MpTQLL+E/Z+TriclkuNMPFm2qjELnodmniQ4Yvdo+oPt
tfISRwf+gXTyZ7j4OntM/+Dzi4XOo7gc2ePzc8N6XHcuadvCYjKC6oQTvY3EWeXc
nYSfOyueEintSIlkTH22RiZuX0P5pnyd1ND8QocfLMaRYUc0++Lq2LaJE2gxL+FU
yzAYsX8i4nd2BEr8xEYW+i+apM53VIJ6HXqYKH5JvqfbMWnbs3p0fCfpscj6qG/z
Ss4AKP40gUIiJ4k5/Ob8GCTqNTlIPQQtlxbka5GX1HKnVFNZJCCenLIGB/O4YJr+
AoSVFeYO0dmvgwxFFuYyCzsA2ZsxCarNxJahqnnSFZ+WYHyYPugUjbg6v7rMSVw0
KLcg7XR79XlszPXzAcElxYkJUq4jq1pKKyB+yGhIU/gbj1oDUkJaGHxmahnjyUWE
Nc5fPGTMkKPCt7hdwad/ZVkDLE6HQ9y8eraG9lIzU6x0LgIUG2uY/cAI2wzNpfot
+jGigZSQfHcCqaJfXSq2/gQhDz4gaQYqyMG4NLyFSP8FcMJn/zHLbg/el3+9L7UB
PxS6E9UJiUTeuAUUEzbQgVBnEhgpnmYWrGFhd205pcUjqCpt/Cx0xkzMnIBSggv5
7Fpd09mDpQePXbx9OA428gDx8auqKrLvKdT0VG2wIrVtX1ju+vhpjgJNhOiUwjOF
rgPBkkWx8XSOIEUR5n8efLuDZ0VSNp0sQE6ARYLKDPh6E0HJX0upKQ6xEzqpevqL
gTw8zIEmWE0pG6KTboQUchxP6s1cf7ML7qHk5W+XCrzogIGAxUWaTKDZNoJ78GyA
M02XR0ZTFnybEAJYQRC8tB9oaHHXRSg+Quu7pfC/v3Moy7rV70Q5c6X1ZPgqejtI
QX4aMfvE3FTD/ZJOUjuSnVqrV6wxVgXDvpiG3dBV97mydxHIVtDa6kUXM4XEhVnm
DnKfu8bpoiC5vaqmojhadIkfGsFvzFF/9vJWflVlECbvxDQ1hASLMg4za6sdRmpt
MQj7btzJmqRdsr+pk1LNmrw/hSkPjW2JK0JrrCTp5uZWSrmOy/7RTz6vaNvfLX0k
6TdhE6rxFZHhv4eE0TWmiZCvtI8MZSOlHdxmY7vXnBAIv5SIt43KaTGI1Q6l5ALY
A6xdXfDt1OsR8vqlmqZhWF8DH9Abb5H+arxrkne4rlaZ5ITUmzbKmT853norRx9e
OO7Gjg3HDg5MNfA+FPcytx29UOGppn+uLBkvHuSgoO/gTMyjgOOavq0saVMZArqD
QcEquiFOdTgzzvEA6pSjZIhFKbiYd0KahiT3p1odBG0o8+7j+Nn25xkH8pl5oOXB
xdTVQKMSP6cPn1GryU6hanj7Ei6E6Gsv1XKtlwNBZKZPY97g3EhEaJ2BaJgGUwLC
cKFnwLD0VObiQbAy46hkVQ0QQy7/Zr33HWNB934dtTyCYczCL+Hf5bEIvKrV/92V
FkieGo33/wIC0ol7ybNLNup9BchvxGty34BLBqgjkdsIZjRiXZhZVIfcQ1bMxPXV
EPu7ytJxG4mM8fF0nDcQpk6EbbWbMuMGpa8RmD/+pBdUy2ttP8Ndi6MAnMow32kV
PJCeBuw+tvneOKQ8ANyUHCA/x77UEW02dmnkFtRBzZASZxKjC2AobDponM5hwRHi
bsDhVVMaRlLnMBV4y+sVmYPUKvBmL9uDsJN+LGRe+BtPBeWP22lPeqp18CGQquRW
6cgyEyudEcFGH4HCkVYpps229DBjARPERkSwolNbr4ccdmdXEcaRNufoL5V/A100
3aQPd4BudKBeSEy5XN+DXjPu27PbVOlf/F/mkrWl/0oh2yI+n0gNI1s5HDj3mdW7
tj+qmaeUyuxBqEET2vY1BgHuJqKXaOMGKE2q51lP16o0g7eSsPNtezLGg9kpc0m4
IPRMvKPfSXRSMPzCb2wfYUId/hNiedL7ZruPnL8yaVgDTY9sw1hJ9hvfW9Qf/snI
m4Gso13VsGNVQvKJySi4FvPVRySqH3WndDi2OaCLFFBFCZQYuIrwMrkPF5l0IoWz
nWezR15NzWvsrs89K+VuDKTPZf/v6LsdQWkXllybvKUahNmzuMlU4L/ia8qaZwkz
nevULmJXhgrgOcD+LtBN5hCIQwXeYEr1Dyr1Ta9TEb3XUGnEPkx5t5exx6vTWj8l
xoETN03aA1q1IhLcBdlUxbZxURxguOpKNDZg5t8R3vFuMvzFxV/A5zVaod/O+pza
8ArKDxnZUqVaoFnrOHmNNgomR8P/jx7jxKKCfL7v0hNjQkXjt9cdb/u2Lyl6FtJJ
E6kyiAWFick6svaPGRDPJQr2m9Fna2AZAj9BvtS3Lu/+kD3pcmlUVlSjXWcOqRTq
PPyq6pn/pI/9RsmoaHvtF9q4zIw1dnIsZh3l9dMd0v7cdpwipRpX81If2kXDHK9s
Pg8f9knnSyifvmf6LXskOl+4Sbg5GbDuWzfcQ/s1Kc5tqBlfShYjJuWOYFF4TGgx
d0f+YCmD0rq1A3NFqwuMDABoya7zKdht2y6jEnedo0nOnCFgJ8Dko5xjhtdom1gk
Shz2pEyndX7rjK0gWRMhMung8kCuI60fF+YIvNn9iOsdPjgLFxXyWTMV6i1ucE5T
df9xw4ktTePy/n9mQh/g5F426FfShs7i1iUzVNK0CoLGbWZhNUnC3f3kZD3beFd+
b+agAmkq2Eurlm1WD4yG4FFf8QZod6Ps8AJOKdWFjPKO9ySKaxRp0Uc/AfdXRcyO
QX9ytUaqOo5KjHe9mxSprpiAHD1X1hk7ywnnXZTvh6ItXTnF3IBnKoK840klUUKC
okff2F3qi88hbY9soZiwORFRsM1lwIUgTkmENj6XPSNN3qgM+RNPwCaqo8Y78RHx
4VsrAgyPi2KyDUi4QjeSz7OryYfjcxGiTGo0oTpE4NZMifKlnqmp+R9jBtFX9NId
2QbkQmf7+I1h0A/i4H2eO9niBWWWa5XWAlszxRWyEgOG41din8rpsQUTytuwmBYb
nJ+nFUU3lelAO8whKDEyUIQAtOh9EguAPMEBiCCO09MXD+ZicSlNoPMf4Jelg18h
Ti5wOylYLzsciMG/E5q8bIa/DfAbwAZTBQh6yUqh8Cdf5tlumhFbRBGuKkWuvd1a
USzcpxquJXgquFSdE1pDlQ8G/fjPSiMZTq/xCf+f/MWwDhF82FYcAzF6lDrUqaTG
94T14Otf3HWB76AojWoxUyRHUyLWbuxRHp6lopyCWIJZayk5lakAAF18Qr0XiXgb
4xFHOepO6JDJTyUVHdVXme+QdHyZDHRsxZiMc6KDPvCMYoMaQZqp0Z8DdDyeEZz7
H2MyKfG3dearozWErA++RQJ/ZJXPe/DqFjrMtvUiWShyzMkqnTOfKuICyRtuQLkg
ivat5kl8Y6EfSg8URAioVic/Akk58f9m86QJ8meKcG8f10sK4MADfVYI7T1+ulBu
YrOGhI/lJ52tJl+TNrIWQUGbr3oDSTLYV8YovP5EvCrh+XJqICMhwnEFfBQm9/l3
2hO7iNPsO3na+BTtxP8NKumrCZk9C6nQyS6EWnzWGPpmJLI2a71HiC01GzhQ/v6u
S3PQS9LPR+PJlai9oZIhrslG1kU6M3omWRQeBIBSXEzIrlFPfDH69mW6uTTqJvTX
wdhq5q/FieWr91gWaR0Vq0RcbPwpYdLVzlxhruA+Grf3edBplXSa/jpds/fkXl3/
V7JLNXpwPaoc0U9UxUClLgY9Gvb4n/BOQdjbMDGNF11pBW+nJ/wNYt2nw4MFz3JP
u9G6Cso2YHlvq2EGu+doXN8pNBWjZuZINAaTKtQCET8X5gPaan+0s6UUZ9hWWHAe
O8Yn7X8WdIs5ehzz+OLUnm1h/Dqahp7tjyOliQCPO8W1/j+Tn6r+rjlOFS3YG3lJ
efCywVaGZr3KEdSUM2UeOy87/3iRfS2YlV5i3Oub3gxwsH2kxwA+/ayVeHbQFQrT
B3OT4dwWW5CuKyJ0IUg0OSpaNtOue++VJG2xdRMWtHIJiOuDkZzjukdZCJWCCgUT
Wu/JSSUswWDG1Q9bJ/iKjD2fy1zKDHSYLK7rUYnH+8i0RHFDYY9HyJrcugsYAiLj
9CNsGAz64PGtGhnrrjNmMPP8ffkIkf1n1cIkR0K5a1UzlV7EqBkWvz4a+Hg3yJ/I
/o/Clm7sky5KT9yhYPw4yM5nr1Ic/NLhUDdGs/aL5qlfRgwsU7CKQC8797VlOQZi
XdjBbkHVBs1wCSJsd2+ib5MSDH8sXoELqFmoexkH49CLPXouUOWDNRFTVib8pUL/
CIIZz/aA9Gvi90wcAOEOoVgvl/GJzSHCBTawfj+l+QjeVuAkjUu6sZXa7qyp0soQ
YEqUUKcghUahlj1aFxznYQWwpwZtU1syLV+NhZyXcXnjWXuwb2l7qbBeqBJr20GP
SvYr93NaEu9fQo7rxc6k7i7JeGfX23VQf2yx1ptN1VETKUxoQ/jwElf+2myr7VcN
Vvw54wLZtEip2ZDcsU/dDoLbENALROyvZAAvWZ/BmYeusb2kerlLU2aibCI/MnYI
cDig1dHbNVVyPN1H8nd7tZgXhgj4HoYsHXwNEjoYgrzMYMOdIPfYNw7mdAf/5HQx
QqZv+apQ6wg/lvNXHIc47ZF3mtkWM7t/tgU6Oth8gf3nl7wL08SXQbNDF65NDJLK
TzIrpZV6UeaJEqNH4l7C7mQU9C1EtBwKnZrQ/IwBI3jZtyfbQgDEcVN4JiA0sxxG
cW7zwMG5Cav8uOhf9gl0TnsWy9xod384ah/5oeF2oGsrO0RIQXsiS2zifCVxaw0K
zdp89vmqvyYZm11hDJD1U/684qVcCkpi2XjzwmeZ+GT0DWJuy4V7yGKRlZYbG1h+
WgmqssSzNqQoAF8FACDVJBgdpzT732IJnpzVcw3rLH5fSAlnnSn5+wE2UO2JaeO4
0TtFJP8YCaS0EDlyWxO0pq5hmI/LVaIEaK0yJYIFvJ8TAqvnRF2QIgDEfcf5sL07
yttowguvXtDGBXsEsP1NMbj06GpSXEQy2NeupSCExxwGyjKgf417qfFFaEVG/pFG
foVycwgvID8oRQ/uMAyMbsxAoDbnhBAsusRd++0ThRP/C1ACoMLAR8Er+0evc78B
SNTzmFJCxHzC5OqwGcx2VaPWN1uNhey7MuLdaylS2Y89HpN3589BsKhUuAH3WGec
PwlkAxeXi+RhkdBMeLvayuazCmMAwW/I2gVAn2czYjh0AMvQ2ogXUS5WgWHPOXH1
6a2x5SVl6+Ty7ye7Lt39vWmQne2Dqd5nZUh4aWWyTr2GgFFpUUYSWyvme1+kwyMG
CcF1IWBmxwfeoAQrik1obQDgZIDPTHJSdKdBFGRCH4qXe4Hi8oREDY6buSEPIKZR
O4MGG97Z1ugw0wKVNBszlnyKkRitVSgBh8SW6U0OIHqKrg5Q/9eqQwn7A7O2Akob
rR7gJep9HDuUVNhEBX5h4UHpLeHWADJ+muInYa6buoQwACO/AEvDTPDD9525ftu3
h4S1ebEUMZ2RRqZ68Rlu2EOEQ+gIGQVhSJVvH8Faw5y9ntu8ryzKdM7G3ge2mqEQ
htIpqYzBo90LQVVPElhZNtiY884mmPOXmJSGFM6CEV76qxlIY8yhXZLXDSMb3rXg
o9DyfY7toy/3y/XdNYAJBjOKRX1qlfARS3MKyZ1jOOqEaVZOr2fh2Q+SzuyAELYh
ari7MC/qWIo1jsRWObY4gygewe9uuO/CiTXy5sztXwfgdIvTQWxFGYOwltx8kZ4u
wEEKPzRPfxhPf0L/GyApAauC5ytiUNaIfcbdpKn/UpY2NuUJtus1ZaB/MuiZEW5s
VuTTybMpuoRzNIf8hinTMwKgBCjP8Mx/aUnR4mmIi9hYSa29LcxLb8F22FETv/hx
lenmP9c73UisnqqestjoC0kFd2JZZJSiSrjnk9ULWaV/043TAvSGwZuKDZqOL/Pj
kZBjegXUZCjrGxvG3UfYuDy0ScjRPUvZNdmt6R0aMD4KPiWsU8PxzlMo6xM7iZB4
FaREkwjbQEQj53+1QIrJkzXH2DJ4IX+7LL6FEV0YDukAJDPEfmSIeXg0WVc6sx6u
AFXqna6+enFiaXQZzT1QeXLAvpO5XoNJAeu16kO6GUz2iGVIcBw15czJdY6Lwh2D
5+CR8829fxMmtULbkHgRl5I5r+Zp1FrUwonRruIq65ZwYj++gLlFqDMN3c2KMyqh
PmHFOfQ0EYa6y0KdJ5tMMGQhWXkp9Krb9tte7q4tSmQQ9edjSO9caFKsPnqIp8UO
FjOc40jJfdM7X6k9HG36/DxeZRxvHX9bEKW+S5T16KdUAd4iw7hkMCcPmx0+gagT
1RmaYBOR9+0IPs3madmGsnQirrsbdfBYVuioCi0bOSd+McV0iYdH0s04M8aNC6Qv
hQyf0sKo4EqdHXt69jg8dtzSUM0P7SrDWF7zFGfZJLQGDrgCQeTAACch1E4Qgwwj
nOljmu7F1VkjZT8ByPUwS+xneTzcnvBazLUXlkAgFGj3M3EKk5hLBqIFv/kYC6PY
DU4Uzxk/pQJs+HtxHAq/oJ3RAhFjzaDBWSN2Uh46rQtcoLLWlG9InqGIOLJJtRjD
AfEwBLe70p+xg2nnE7V3Ct6l3CWA+fCdMgCVLUYaFbOkcFHAmz4swEPkCuXD9uXV
RHSF0wPy10PEUywiUYoGQX2NRo4rMiF+MJag3QxjOVZBx/VLMfaxMo4YDW+Q0g1Q
plNscqoZ6nlkInS8s825dYJVUQAYsW0CSjGqog9KRmrjBuKtJhxvCX6bmyep++w5
9NRqH2vR5wzaw//+HKWXR/uGg4E92R3sLh39hPV2ld9G13NIGVpo4dn9kIHyLniB
Cn2vJOpc2Fpdt+o1qZ3xkfCpDSYFnBm6nP+XfnvFQ60BKjE/Kqfr+l4nGXVycd1d
pcd2QrBpBeA/iXNoYugkJ2RZtws4+QYc136DU5XZt+f1L28MwWYJbLFjU+R+dHx3
AS2UAwdZU7w9rShwsy0vCy/RgPaQkbZll6jg0Doz/RYxwqxbaGIq2vHQrAKHedhN
+tVGVHzA0VaHv7q7C9yaTChMwpgD+xxt9QyqTGYvFG6NCD/tSdd/SRqH34IdWkor
fwR912ARvhCjiUb4p6In+TwK+/sFElrdkc5wwhGam/uAZnrSNtlPorrC7J64KhO+
Ab2OFFkx+UUv0BQ8T33ES4CFpSGX6py2EVZgHbmOCbd2OAXjdlLEqTnjswyGn9/d
ca9JMxe1/Zdzjz5UKUKW/YgBN3IYtu1lvblZOCN8hTmcmvmolSlVRHGZPdpY0jsN
2nwfL7m665hCmbSYhjVx0sIGIPxM62RSer0KNV73/VDe+TNf3f28D+TJ223XUGfc
vDcpMPbNKdvf7sUF6gOQs+ngAvSwKWIavBhS1JGIrFLMeez9j/fSPz0JAeyrEbFO
Un3qx51loofwkQTxvhLPtRRNJ73fEJ9WDAe5mh7xW3fZ9P43a68rkQtgtK7Y+A1Q
GdduS0shgPgJfEMWkx9wsiWtWG1lLaZr4JKLdNpI71f2QfwMpwL7YQzjo1lbt7Dp
zqrbjlq7W6hHbumZEf7C/vtx2rl+Zweti6PtlBoxbjAXUPDEkHboIkAolnOgDkPt
b6BKlwPZhRg+bbKxMeI+QuiPtOwCC02MwmiXvlxWA392cml+p0ciQb4R3Vqm2uDQ
qWx79iomat7NzhbRlARmstzkKMi2N0cVeQeIqERO/QHecucc1d9qWoPml7cQoBYK
mojB17bCMYxWn8P84RQjJH3JZddg2JiX7FQiwrh/aOY4grtTOx2pWDCnbThK6hLL
fvs6V5ENhktDJTMxws1ASDfXyeieeZ60Jcmr50iZTUF4aw394Y7tl5TbNU7IV97+
RaT889NNdhvUAZ8cHG+EUGiTjRaEDiGoR15jLlncXyRI6HB9SirA/MVEozzO3fiz
WUDKGhAiVCMTAgtuik2wGjIjd84gBhGCj6KlRHbtENiAcgjnmU/ZvRgpLfuskP+w
KeQOaQWOh1a5JaesvK+B3INRfO4ha90cjiMCnsaL6PPOO0JQYhOkcv+DX3CYGoRE
PegkUdQNsQAz3pKZD/jpZIdFsTV83bX4o5+sEBiaSh13crW/ZtKJfpBCcRrNvqdw
DmJrbth60m7AKzjcCf889b4wuSbYES4h8m8J1Kor5Tm/tvPQquk/3hmoVQVkY0kP
0MobHGqEdyvamEoIOZiQ1oEMK0V7R393KjcuZS+xohQLdFQfe5rx5eGtF/mdBqGV
r6VVeb5wgsYoW7DLm4HFJBFA0ghdL7UzKjEWHGZW9JA3pbJK42Jl4t7nsWcu31O4
001Ma8xIIb8UnGObajnCV+el2mS6MxSdD9cG+7TVUP3K4XfKv0mKJ4Lg34/EsBq/
EwNBRewbas2VX/i9fNm63vorBjl/h10Bhu/h7FK9V8BJ3Z5gWKHstl0oysNzXvsx
voFQkV0EN+u0xS0twSwSTJq/Ftmf6ih3z3qnCdykizS1WcH+pETswx0VGUU+yrL9
Xv+ien3LtteD8Rkf+ofa7ZEachbwuQOgDp8lIUkpra8aU7cfwxDbtnYpMiFMJE0u
Txfms4okKx23r5E4rp8oBpYyn+wGOR7KYbfQeL9Mj28zkOdd8cEmSv2T+h1L5RR3
xHW7CM7Ntk7VYDsaTlcf76MxMKrZU7arozjTGaTyw+BSjhwnucxO0fba2TNJInum
Mw9yrVPqa0Hy+QDJEMALzrkb3VjUTJfwss5/Qm0taCxJsj2iaTM0ekl47NLw9o0A
egvV+st1CD6CoLqZH3RC6L40vDc9OysJ8vJVO85YeFSFEjvdnIUeJlEQg1Zq2HS8
ic+C/KLoQyl0MsCXn4wSBIUcVABY27yAyU0QzkEcGxdUR5+moMhtfOlif4icewFc
cMg/dsBJkXILEm507taqprsCcy2xoUZnVcpGVQkB+Q4r5o+Br+Dz28+7i0DmoY/P
ClISHwtUC0T1VzT01WmDyNKZ488X+35WrORR1DeAVRCG8ya5DPp1UbREIZwdhHke
JRYSPa2kPbrUZlqfuaRjYvLFVD3FcCZ4tgP5aapd7kBTvtQt8qw3nn6AGK77RJ9q
Y9nNpid/LLFAFdPAybSbltIlWneEik5AAUCzO1w06xFqmaCtdu1l7PsnuOOvD2Il
q0MXpz67USUrWyfjGQJfA4T6qv4ejbby07cjThVIButFVgngogIVht1HmHvT20sV
b+ponQJgpZ5CV5Rht/6DHLUl0duJJEy5ZTSJAY1UnJfG0azZECdVamUBEJPY9tZc
5FZU0or5JJkKZeJaW6VNbjyWFJaVYW44HwMvgp5o6jkpUQVDKcBbQSh/DE2UmIJ/
AWeHCTNfC11JapB8wK/TQF9nczpy+pqGQ8akI8fl/l3JG8EX1ZCkvWgK0WFuWTpG
zSXCRfKrDZS4rXSUDD5tQNoyr9/oepXmMXF6yQjz/j39G/sk2rWkkKUsm/hbQsU6
BiV0ySHQ22BsPLprreBz2rQyiXD3jsDo9gdKE3GEQgwCo4za2ou4hbblk4rv3ITL
faCrSSmRpj07d0HAebNZcZG00ZF1ncZum/Ep9hptGbHXJ+sfTa+FAiMuxHpmId12
cHSZrs83wf8zH9GKPvdI25HWI4MDmXBlCBZLaeZXZVXJigJLjA9M5bjG0a5MVW/a
nAW3ODPzLu863WAkkoap/uyAgkMhkWHVyMXbb25tenvv2yaVyorZXM185fAF1g3B
VMsmyViPIaDz9EMhWwDQRBzOKzIlth0cP/lEyYaByL993AW079YS7nyZGgAWikEA
IMDlG49b5Wkglh3JE3h0zFW74obe3PqomWgcqwdp7Eo92xsbPQl47v7YTNh4XAwC
L704/1Cl/wvrV4q9ZStXJhsmOazfisTHGlBQgv7Lnnr9qdNAM2x7pl2p1az0Z0H0
ik/xcB1usvK0zp0wA4g+WY0Yeq7k2QMIzsEBkESKhZjdS1uhrFg0C5CMzoltJFYE
0q/lOJi0telqwcHgrtpRWspjqydh7P22a+clCkjzlBNjwTDzuv3SPoikLMs0L27M
dAFjfNopRtxR11K4uUAcl2p26OY2sKznB3BhrjavMCv9ZG9hyqZ5kuBGFGb+p6He
4Gu8jVMDF8G2Pjrnu9lQrE428nAfalUk1HnPXCcb2vkGn7xfd1h3Dnmgogu7eRnJ
wYLzk/c8F0z0tnJdRiV3qaa/rXRT6cKbUrmMHxCYutfI5MgPiTjZnsrDU5ZLIy+I
5/N/Y1XYSdE7rmFz2xMP24JPhQ2XhJBxclIkp2ph8jWfXZ+edZ0wDXCGyLJhfAQy
hZo2sWf2RhTT5EJUk76CvFW2YAhZ6tBXS6SAwpZTKyHUv5cVE2WipIwA3xD0ucII
WIkx36F31+BJYHeYzlHzVRPRrbkWiRJhf0aua/2c04BTGzhf3HEbeejnxiS3mnDV
/wh/AEd66wMD13CvIczGd0bSQFVUoYdNRBW5zJcYSb6eJfincMsA8n+AuZG9Kj3A
oAv7a5snE17wSCk25+qLDYoCoi1CIXvL7cs6PcbK84+LDYMT0mmsaLh70IY9udzi
luot2+HZ6TvdIUiRddz+tfpfI+CZyYG0KxizAY4nNWaB2VLg8qEUmZCFlEHh244n
DyUAqhCM7kuwxtAKUEOMrqm7aJuZBDo9R6QBQtO/yP1bVhbwDX7+/skXkW9HSYI1
z6qDyu+81tECMjJYMdDNh8M0d/UtWQYhvi5qFq9oDLXG/d33IVrHpdkVwKuQM+td
kkcm7OKggDd9yTnNtQpJcbgWm8MVlwgYbZ3n0W1TMeLg6rhJI+ck3lHdtqPgvwYk
lQYbmsZbDA9d9KpoCfmjB4w7e0Ag3Somn5VYfLDQk+2nwJY6WefqDHhL5Usiwq67
yPzKYKe5pWJiGT++qqbVxBEAMZFIvpcp3rXm9RginwKR1Pp4ej3aYBinojv4USZT
Hi8dZwnk4v+34amoIDyIuZ1NgkafwPQ93sQWaHuYAS/97Ln+Xp+/dhgv5Ad2JEUO
9lByCQ1CGKe2m3DjyqLTRt22mmx8n/ac6V/LZEOVMLfvkvbNTKGcIy1W8EXuj77w
KNZovm5MZn+3p54cexLCC5nnEXjd4sHCjZZ3EbgxnvjS81rBWa6dImjtKBk415gP
b+s7vQhhUqiiIR8XWeryQMLiIysPqDJz56Mz+fUpQlkSQtX0sCXMpPh9jacwvOhb
iQK5xMOdqyFBacjT1Z3pcMo4mbEyuBYlbuoqIPqkcSYN1iXWJwf1nRKLCwMZrG+1
Gcp9dD/FYxZNc4dt8xUDAqJDrdXcK1ZbM3IOJ1uGL+TCcCIF0jEf0jSNzpOxZ1e/
4rhuDT0EOcg9MWXWSYrEJ3Lqa65naZH3Osz4F3Z9gHdR5NyXGvn2ErXVQaFLr3aL
yv+T76aC3zVDr+8ceO4qvIfWZJGbkW4tl4RQhwDjFRV9y4O82Em8fwHbQ8zv7HUO
BKnHYcSX00eMh22EESskvwPjN/hJHvs4lkaDiUYTwIfiE9L/EGlbyJHlxSL41vCw
QzT/GH4VvVnsoe1mVCmitw+cVXQY2iHpzwFV8j9ouj34n+OMCnF3spaL9gv05Xvu
/zx6nvvlSmb47UZNARVF1EOpobY58w/fQIFU9yXsc2PTFckIqgLXCRP280wRrkPt
Sk9V+MC+/UTfFSstonCqt1ov0TPEDMkIdRYE3eHEo1HCfMO1PQg5jsh2Xd3C1iGS
4xmyK7b0hpGzEEHqFi3dJEa5VqTOLeLScxsfzeEwch6pLZgx7oKgzfdW7JX4B/uE
ScMnIX43s/vZlGu3d17jHV5fL17BRGk1IBdZmlzZ9SIyYf0vjT7skgU0QRwhMBsR
tSfIwWgsBhpOoPkAb00T6hnl4ku//mu3nLxjbmSNdjohwha3Q//aTOy77exyYE7T
KEJgmg/H5cRjh/pjcVhXvgMYo/RAcBNAHTwJsYtnCj6TItfu3IhHA18ASCa3lSvm
fxV16GW6qf/eHGFXzpaK2qlDKIZF81QCx8KkM1S7+AgqtNzCvzHkNxJdZrquKUV5
Z0HtQl+hxlXwD38lVlOmTdEwOBbLQ8HpXvj/Gnp5Mx4Tr8f4E4Imc7E3HsPCiUZ0
Ou6zvKXHy15e6IAeAxgyj4KFIZ0yREY/a1HotCVFSQ+sqp7JEhbmry5NU8DsXbnx
FB1tNJ6Orx8YrNzK616CPqdlyp2A/MEGW0HK2rRVjhvH7R+WRI90FVaB4P2zCI7G
4rRrCqGgUJ0oHYgQCtd5mF7eXodu1IM7q16nsUzl/ow/zxWdI1MgWyIfjhD+BmgP
+XpiqGQjR9WM7oO8vYNtFPro0Aqne8fUjgYS81ixjtr1GZuT4v7ismhNVsOlnvzg
MCVOP2L6T4Qd7NKP5+Djyisv+WBpbYC1mXxrX1egSAuMHd4XIRRiI1pyY+FmdwCF
hyoGqxOHe3uu8JIaeiXLU9suRzdi/6gABn1WmGvAAPjXgE1Xt/g6Zi3NjKNi/0eE
X4YsGv0KRjhLQD3AKqkuDmdBhBVRLZ8LE5I9DfKYi13BlYh8aIqgXYKsxte+0Qkx
oHh187yqoGwN0xEbPIFijVQO4mQQuEQOCAMY4f4zPsLN00y9Yj4D/xMGsuwetN2c
24lMmPHw83SzFQsOAf6oE4fCgIZZOJ/qoL2IwNOJcc0VBqB/OiZiUSUX08Ba0aFw
i9lPkNYMYKM7ApOXT2kJXjT5aTwhES6QFK3xmTGh2U5gxjIF6NI21QiXLExfVRBO
lQGClT4gZ0tuDbjyr1hCq0GbCjGN1jOV6EeQcQDSuLc30YZvpKSFS5jqygfoiN6t
7hjxD51Egl8aZgavuLhuCX5u5mTMDfIsihDY+lteFYy8eFy2rPUHvqZ2rbFQKGSa
QAgfwjt3aGq2H4JirMBNHJDeEpQFxxfKpZ6UaifqpUI4VJ1uwN9FNfe6VCrPNjN2
k7qM+Nc1brteXhDWV42coBIWqzngJRy6VnjqfwU6G/V+Snjmgl7fIhpEOylz/Tib
4llfHyJ0zJHAm3b+9sb1pc9JZqSdAX5XL0OghE5H5MTPEYSgt53b0vJg6L97bTZG
moBDwcalHtAnD0AsmJgMEwCZwpRS5D8cgi26AQFcbZqdOFD+6QrXiCijTt+zU87I
FrjyCQUJ4zRCjQIGPZAmjKqshAoORdJ8Jl08yEl7VtLZL+NCsmZsDadYLwdWVkRZ
6l3KJBtw8H+6ZBo4qhJWMzVgm2HjCaCAdoZsPmj9fsnz65vNHX6EjeTkSegTsIcp
czvEr7kc/RFULgnxzgnRMtoKj+oZe0Jzd0ztCSxnU3ChbxQrpEJQk1d4Seb/jITQ
o1SRGRWlC7TycQvSBpIKReI0CDfVNGm79U6xaPWJbaO0wqd4dl8Xabt6zMgRB4Fq
Ox/9sUynxIXwKMMpzxcqMX1MHVZdKoLoJqx8sJalCU4pcudepjT1e8orGUZnyw3u
J0+PWVjwk4X4vPxIbIEMtFvv7+fFtDzpNofeq1IBQ2UiRyd0Kj1L9JNuMRQu7IiJ
+MkVZKKNhzAayoqeW4lkPLUEpL01gcsXF/T5JTtmZnDcJsCatKbqght04kxTyz9Q
834oChw64ZRGdOxcwUmoMWMpCxIFGzgWUNPu1RNcFA7VUKi66HLy8cwqjOIpwngG
y8dcf/g9NEmlgXQtQwFPoL20SRJByX6WBRAeEn/OzsbP6ZsMXOlm3qdwVmKXMkFc
wvM8Q1lXJNoKYi06Wzh4WoOi8mpfmZM/DjZHJPtNkPVEspd6uvNSrplOPZJ4I36i
ZIhxZ5SGMDMQp+ua2zR21RO9LOI5EAn/iovzdlAKbO7Fz5wR7xUjucbwlPfsli6N
D6Nk/fRbYJpY9vd0NBihlwOXgpWhXKpFyDU+0SJvuzdgtVZKBM04CUdO9Oc1v8Q+
kd1+Az9dBnLT+ZjiuEY2YBWPLis7UeF04VZ0hnyT6MWT0VcPLxgsEwwO9VPNyVH/
vC2fxzMD0dqFZw+0UE2OpTVtumN10FIULqICU0x3oBl8VTzyP03AzisJSfF4xbLi
1sEDKiWU1dtXHPpt4G4CcDeKqGq6ihpqpwAWWvvzTiS300DEhLxXRACGNOUGEH20
M2IMuUTIapARYaPLpxjZcb0ZHIcpPFtlLvGa6jhBVw57glwCIGViTJ9EajGm8XSJ
GIje/AOEYqzqQzdX2oWCXR3lx6JmQHY1UyxCJuf1vVX/bYhem2QwnRvRwezoWBK2
iTItHFp5dfEWNePU2AECPhZdoUUtDx4KmukLbgtLEEbZWKcF1Q6Jdyq7xbRB26eJ
BsS7bSrMvqjzi0gZzbUeNNrJyneWvjgqV9YvfVWM2rHpYRruIjLv/HfPsODqGBBi
R8Ij40dcN/2KdZyqVS3b4ZwX8aSn5QdaSDng7YF1K5ACACY47fEly/bhFb4/eNtM
94MSan4VLLrFHz1makWU6XS7dqYR/eAcTZMfLKhugDciJl62mQcn6Mox5i4DaxE3
srsuu1l6YF+1xsdCBuMPD1TzMkyCeFlROjdZLaUvYGGqeGjPum5EchwDn5/reoRY
As0K4WxKITImiYZm8++OV8qAiVhvJRJhLRrnPKYaFmbFLR6qiG1rTMJGpIivaVkZ
fLwI8swHsmPCgMzdDUrnRrUNHTAv7NJPOUq/LnRaPDNx+nKRL4QzeUx4Bk4Mrm2d
q/Fp3RI64UxJUS7c7qtYTwpK7bkmK5jytYeF0C3jm5OO7e1Kz5zcKPkg4q0QTtrf
qxJGGB4rJNbg+uYX+pT4Y7FUD1NPY6w1zYYZRq793S91nal8wQUbcQ4lCky+ZNu5
afd0ftOkIBZ1Hf8jLsDW6HawNr4AK0xCXeWcbfCECosWii50BL1Zqr+SsCS8lqNj
1TUQXk/q0QHWbl3NCyQltgRv076N5Y26kMmxTfgVd+9xxXND4nONhkmW3ELZ8z4U
w5b1vl7os42L85ktSCm8OoNUWIHssVjVzPVKn2bg2Z3HQQyJSk/ZZ2oEkvGnZJk+
MIk6JyJZcVCGuZkO5n2BZ9zhEC3TNXlRGkEQt44z5l5zCnwThypgeX6HSSB0Fg81
UqmmjURcWU2mLSCnBVlutmMMD7NS63HqUCjA9FTqQuV2X6//iupjw/J+Pb33awdS
+1+0vza0PCcwPah+OYc/qOHDT29fupEsXCO/inCOdy0T+C/MZaHcxWOzZQL6yCpg
1TvrpVsCcqLGm4NBYP+1uPGvUQcztty1u/4OyrtWWTegH/X3ZabPn03QJ2loDGQT
1NCOZRo1700PKyrNqN0thRnrfEqOJQ2+fvBac9HlXwzJfMmbUdPx+/8puZIggsP7
VjssOsa7AASP9jJAN6PVB/OIDxOzGolOJhBhqsexM2dgIQvI4WWozt5Pa90zmWQd
aymA+wH0mWZidjtlD+9FraPoASj4KYE9XKIhhSMQm38f+LPTM1M2AA7NXNLVB5wa
lDlyPFRyFiTt0/VZJrYPYxZwHdYgpol/2TfrinCMLI2h1sMroM/aU5rbqYi2qqav
ULfoVTlfCJieQ0soi/5cS6Y/OMQDHlWrs8WBIcoCh6zs5yAIz1GdvkovoBO/wxXt
DuYxwcHquRtoo/LPuBEugMwcf54v+d6PyT2qqH7+/Lg6YZz9qRaxUzZbF6aGatiX
uKZRXFYFPfC1l6uNalHLBBRyts6UP76X/h2QSt8A4QsOqC0Nyf4fTYN32gkwejKM
LlXkbQRKG3T6imWAypyF92jXJvM2dT7cTxyqY7hAdiiOi6PdxRVIlvyzcPx6wRBp
34ymKbiAYDu/uJjJ+QAgh7D/JvASdFqUK8DGjEq+RVcDEIn7w/tiqHWqwzD51O4d
bUjYR+9vZZfOnS5idH1P3ZS+iL1ZVaK16kaA9aKeJavAfAJEIpeMOA7OIy7KN/Ep
n+HN/YQ8CE/6m+iO5YWO5Hysnbz5HjMJS9GSXBEpXk9BU+AN1shR81FdUDwwpHjb
uNiwWnldPefCNMm7rE1wW2eimZR5EFoHh3wXw0M3hPQgKGSidy37/8ehE6JvryQf
9aWq+4ceAAkWx4m1jUW/Vp9UrEmPIUi89ihrExqseaA22nttspcPm7NRcOdWIFPJ
85PWpckqrm7eO+bKFhT72yeSe+7BncFYiRKeeyhu7zuT4s00c2YDatvUfMWSYfPt
6hTA20L+L9MdH+opLhN8cBdvutHQQTngVoifgLzyERoWKm/TQ9lONEx6+iOufqoz
+3bYw5u4Wt0C7hUPNAc5cJuD5SzzOGpV67XZnTSFHI0HZhvWGAHI+n8+HnR4i9XU
Gf1kE6ogoc0/MVOVeRsNHgYkMuesSPvmOUJxNzA/mtbQqpmXkvHFn7HTgi0aofq8
7f9yBbTzsgonP1jiyIgAm36QhWEpu343eTttoSgGPr4mu3y9gsIYAqTz9UnnDiLO
KKs/w6XV4h0/uaZSnvDWmeOJx9SqOYYNnonFZ+NfVgSdVjpcYg0eL21Z8lmNG6xu
MBUUc5pNKsVZx1ycWnRjouMMJ2LuO7EM9VmMgwz+dtLEGVpwHWYzBrb1c76jFg97
8dgfNYKDfcckCW8bx3XIOF5UGUNkC1ZsPKBeviCoRX3CmBH2kB3Kt5wJ8jZtyn2o
2BfgsMzG6kHDwVPBjn3x/95pzwT9BTjTdc6y+aFQ+ThZxINhdhaYsdWupOpqMIqM
dF682F9w3/8mtVdnQGI0qIGFnSfADOdEIeBxIe+s/rmwY/SbXfx/5KOhKU5QyR8n
a3fhRGP5KgCJXw9oRsnLYBE0RvX1KQzpXaI4ZGDgXOnjcNSR6ki6MRfQ6f/3+xMw
FES/gnsSSbEk6TmWDymZ33SSwH8SMbKFfC7mXtvornHy8i2eLfKq4q2ohp6ZKk3e
LVujJ08c01HrnPzEVXdlGGZJfxwE0lViQYesiNq2YdGm49w+6YuQOXRjEuE9JXQH
gt65X64IfvcIUCGWaC5bT/7g/T6A/jK+4ToX4cd7PiaUA7AsTbHTrm2KvdcEISde
KNoA8dqt7/F474wgkQ1xXMgn+DbULv1YhuDn0erX3y2TVJjldku3T/ZRceUB2xu7
v4/NyIqDdaq7lxqO1bsoPUr0ABDk8ClS/GxZ9TBTYMmr7pnoJqqiWLfhc9DWYl4w
jk62PHJ5l+KzAESseLU3SjZ2Tjz3MUBzNKv56Blat0m4YVZrhTQvGQpEbYfbjaZG
xSN7sxdS1PHSQh1nrg1O+xomLw8rBrB70/Q5FjK21RC908aUQHA6VQtHdB0Gdk8P
RrTHJ/k2HhkyseN+nENV72MMjP64stloNzvbQWoZhWpKjoMByOXAR9WjnSUi/5g5
L8a25lzDCVjenek3hHdCv8B++InhkTeT+FS3Chs9mltog0w4OuAM9S0ssbaO/a6a
43dXBhi8JdBfz1KNkYA15I19o7MPtzgiXOT8Gv3UhLRXvRdlGazo/OtMTd0C/zmV
Vx80zbNGX08Q042jwx7AyRy3z1zVtGrE94Ficbm7ZHhBrTFXSWMQaagpfNeFGwYs
fTpvrGih+zKoQ32OQ7lPgXXXlZDl8gqVvkeUeqKhoJR+YrpxF+PKyMjyXoSRBX2a
f5n/ErZCCq16wQ/fgSrjNdcl15L9rm7EaVIDdi1MVP1d0X61d4JHj5BiBrX/6w50
KzkSg+s7z5d5g+ilOyyNt0jQVG7lMWUQQpjdeypwk7mKAgRF0fXo8C40ttRzmmOf
RzmsUEO1pHMhcicPuz9XCw5grbsblEjwMmEgq7Z5AX13WeblBdcdqIs97iz1WOFq
rYVOg6Nvnz2GSY/ns4ziyxwm5BHrJP4MgOURFrFvZfKGdVVq7hAq1cFESLnzj/NE
BPEnD3/QruoiuvUCXWBcFQUSwiy39fdyTxpaaijKV01kJRStbz51pysokg3XSyB0
R3+/g1wwYqBfA3ErnGheY2tT/0xDgLcZQvWxALGF/YErnu0gTLZrqN3vXhDHNrsX
sTLfIu+ebM6dguJNhnturfsk9hjqSQ2ZMaeiDdaqIA5OY93pURzPQMWjBqQCpqHV
Ks4jUOc+LM6ZICf7BCzbpasX9PMSKU9w9YJHqGLHrTyxRPuVqipPnyyFYFkzJZdq
Pmi51Q4IiuZXbhayaJhupZL+UMjwzy9m37gnTEeECOI+vwNnvbpx8pGseMDKTL90
Hj4TU8Nvv2ZJq86ny+lHxQu6MgjIi+YnPBza8R6VW6xWoIXCF/Kp87vlbv50WIWw
ktF3CA5Z5S9U7cLt0k5vtVXFlJsuKkNx8caxOYjZ7iya1LV7GRBElSEVuINDlYso
YWRH5M+kUjw8gSUbBNkrWMii/5Yr/LimTQjaM8z+YNLtAI0E9rbXrl6hPY+OFeaF
FvHd7/40dVElu7HmDmMVpiuvIMFpOXPH8XHFsetPPekOGf4Jlj4HezGkaiC66WHb
JE6tjq/ZM5VPSweaK940Ttp1/BeY7v6u0NxqhsSD1wMR7M3ke4wGwJ7+j9Hh1GEV
uF8zPzOooorlmgCaP73KvGnMRLhMJzRHa2514xeTrja7XC9UKWtnJ/u4DAsYcoum
gVYuxsOSJ393cvAeDe1rmBqT54scp/gTyA+/E0YZi+wtG9YyrGa6UXF/KdSLhEnV
pLjfOnXp+QdG4aphMpd4C9OgV2QE4L+ApJeME3BqW5Qk+awXQOQNJizV6g0K6rMI
OOupJgDNiyyxfTmvVH6lwj25qqVNbdQAbT28Y3UPIZ87uyo15YFkefDGl8kJAk6X
wikBT7/yjur5sgoCid+jMRYPHK08iEMqqXLoIHFNspoBBaXA2DRDdjDtphuWYGyq
ToPHjiefqzIeAS9Sp21hmNhTci50hQSROEO3ObwPoW5HZsGAMUSCff17h62wfmKe
Xsd1Wh6G5bPRvGVTgenVlnJrSBvjRK2CEvnZiYvOC9+kQulTvoKGVKzq3xWFT3mY
LWyJL52HsIdWC68LB7y1Ilmj0GkNdK2RCU6jv4CCOIihzpyx8r/Va1W2SLNvEkV1
6S7CE4OeJ+CsVd/c6MP9I9nj0kEgifTblESRAi4YtILxOPvYua0bzx0EYYycVPT8
2GVeYu98aBEA+2bT/Ji6ofhjpMMUAfteQpv7rKM4+u0Zuq4rz39wcWM9c5FQYvzu
pqPNqI17qaDRCybR83kmmTSd4o4caxKHbIPqEtUL1IOhJWSUkYvFURDN+hxo1oXQ
gnIcrZ5s4a5uhxhMZZC+mixSbiE5TQtZjQNM74vefyRaoZENGGMmed9sb1h7l3YN
SF/q7DNC5zcG7tSpC+KBSwKysMuvMMDOq5XcJyxj+/2w1VfqrF/mqFckKF9/LEMY
tDPFVyMzcFCfkMmBgH1hQpTsXzLg+jRkihuEHlGLCfRslZtUrKYxeM0vd2En5hwT
3SN4g++L9pBjfqfON3McsAKPUanTQktDDWfg+58sTCAAGNG0ULYzvRIk9JLMtJ23
jGUP/OS3entCD6e5vlebk+eWq0v679gv/qCRHaZR8mSAN66ypFjbHlgS6i6hzZKT
1A2GwcqUPJeUzliRupdz13RUhqnKZOmd7Aa+nVrdnKmpFt9xRr/v6Nj1d05SVZGi
Bnqhubo3CasE8oz8Teq/5eFx7nzqmo70db2m6dfYbyDT67Ahz31G594g1cbpQsbR
qVOpc1fdn+ZjPhpnj7q0Xbpbn4+s3u8FYm4KlYg232b8lnVoFk7iCeM4wmGm8RQi
cclQ7DDnoiLWTsvegjJfh5AgSUUCwENHqAETUNCrvPogN+v8h038liMT77FSQBBD
TQvFxbV515301BGlD2xgI0eXV03G+UcBI3xTy3NSr1KRRZiUd9nXXaQZPqC6EqEB
3W94KzootCxnhVjkb9ssA7pJPR8Z5XLYrCyaRkZFoOHvK4mYLo6WDf7ft2tLpyeT
2yRzjXbZVN18IKCud4+P1fKE7pGvKJv/Q/2Ap9EbTV0TshSC/931xk7jmRLmORFX
gf0B18DQcTLtgqG4Cye4mQbrQltEc7vGyrEpL1LZ4TCYMpMQiHqYMrKIhB63lkyJ
O0W0DKKTiWrJ4XCsG+ibJEyVWnFVYvVjT7TVOL4fV3Mko98QJ7czroCFQMXvdIjc
55XLkS40qPNdhFRaGG1pwUxQ+LGxPXa+fPInJGFBGnYO3bO0zua7DNuYRmXUKu86
6EYAae1nsbwhzRPQOMGGduaVRiMdpj5+qpx/HdQnYicnVLpgiX23Psu/CTDLUf5T
dLMg+UxXoQoB3ZBbdps8rqMHGb0BI2t9GN1SY4qylylr7QdrqGQlMnhmC5ZCoyFb
oOZMRDGpaetwcK54W2yVIvgofmC1xerJvBEhlpupgLB3/TOY/ihTHJfFvEESrWqf
nQ65e+zYHZiKkPHbw++pc2s2wDJhMHdy+lOYXKtiCOKly6UbZAaZfyi+DGf9gh9f
HYnw72WC0REjmxSpl5JF6/HVMOQd/LMj0tnO8W5auXUbYR5cT7ytiHR4hWgzIfty
kUDuRmheKhdLWPPKFtm0LdDHiEo03HCPjHF6pGD0WSDUOd+qTCNF9Pz55NhVjlxI
g9xuXOtXtzQqJtW3MlHe/wzdiDClX1d86b4LOvEI1yK1nrnSXo0f6/l5onqx2iD+
NaZIF3D3w6JG2vdyxb7HhRAOtzIxKgKDd/W3emEutHKnbP8i5P18Ksr/gzDB5Y5W
8ZSwNN2dI3aTrMgYjfha2YqHhqtkvLZfdfF2rFPb+XzAdKxi5eSgBXBvRPqWi+zK
/EBjl0tzkjAIqVEy7x75yx0fUUFKSlZNeEVYKOR89Hris+aVFk8/JjNmsuQ42jL5
8qcKctWnBnup01bVPe+g31cMc6PgudFV2kK1QsjHsKT0Y/gbBHxAf9w1FG2gCErJ
NigOyTFgE/m6kJPkFmSDS3xlNEKrSTkthEQ+kzdSlyUDTUDHwDurw/8keHC7YJg/
g4GEjUKgV7rCS48k5OOW21NY+2KFWMAd0qhHTCgahsmMsloGr5uhVDD0sh5FjzTh
pn5fGQ8F3+ObQ44Q+oeiXUHPJmtJjUgL9Jkisk4EJvwUru+iCOTeNAfF3wOrbEj5
x4zGcRQokmzUE2FiPk17rsHhfHqKe38YVig9rUqXFNu/YICZg/BmnCR9Qzvx73ZY
ZtLJV4wn5PzcT5wGjx/Wro/UEmt7e+IFal9/DiYz5kRU3yGDxw67VQrdjXYUif5l
inMDmtc9Rj6zPXDeVZDZWlWfqXvp5On9NDPjIJ4pdP+LswJg+9bYTf2gobty6iiH
3pGgsfcw4Q6vXHFZayrps0DMuzaDra0ePXu2bFxIV4zCJec51crQEFgmLlRXZ+WE
94ISwpH0Aze91xSvXpAkCzW6JLWN05oDAdUEdug9RcwhSpg9itMkkdoNTPWZU0T6
JIG2I6KMZbUn2biKNYMOmNJp0fx56TZQGyBpeoWK4DFldz02Aa8OZyUsdIV7ta+l
CGwVpLnek+b6VzQ8Ndzqgy+EmLL+B6Kxd9JCQ6rOb6MKBln/T71TnkMLjIhNrev3
baxjQCDfUM231k3nmAj429sMGS4YsqY7l1AYDwSIjtWww/ii8xsZrzbjWruB6MHQ
xau4l4BmoVlGTXX/I9ktRdHoRdHKRtBVr7s/nYTCP6bt8E2aA+chfJFo4QAqW+/H
THLwdeYxy9YF4CNHxm7ZdEwIr4MNC+Xr6s7iduCW2X4Jz4Yi/XqxVLVVEsunUwyu
tsFjisUC+TrgXGA7R1J/eJuT/St7IFG/DH2FDI++RZV15VdPUoJDta/83pUh5HRk
yHOyLh74KslfOockosC9jktspLo3K/n2Vosnd02d+a6ohT379hqSQZELIRtbdC8y
iGWElujJNDccFF0K9KUFujKN2dz7M6I8IMWmM78QUaqDiLUMCclOXdqogVymHsS1
GEoSqrBO7lPWGDEfbTXfppi4B54sujsA7ipqtwy9/J6RDe4KMdTmooQDdfoTygYs
ly+vG3U+K+6Y7Uqd7E25gjZlhS6xzt2raB5R8vyRHu8m7xDzRXoyoaluDyFi3cwN
Kzq2OI24QdAP/tNK2sQ0x357tGHTZZc3Gssl/tPVFbbtexKXBKJCmk5QsPFB6gRM
sU0j3V3Sa6q+fiEkoxX1O8Fi910UZoPI/y6yDvMCzhxhnvTcMZiikQ+C+mqQ+tvm
ri8hkvtt+Ot97oWhiJOyTbRlsaf8u5QopRqTJ/7Ay4489vSVKoiWjw3OKJL3/l7j
H9VWy4+XoRWGUXSwZMyfSjeFB3Yi0EASXbvy69nV7BNHNR82wCXHpbwgqihrjYX6
Wnc6+lnkybGr6pMYRgMKxbAuTIK3x3qC83oPh98S+IAlM38CASsx5K9Rc2Br4HS8
2qJtrjYT+euNWbS5WaerXsl/G3BdrVSb3+JpZt8krPCqXUJh8Fwa6KxXi4XT9ael
bpfX+9/dG8M7IFmJv7yORitZLfswBkSsL1cqjb/k/8rDfRLp7jmEI+VLCpHge7nB
G3Wa38RGDDXq3+z4LRDdAMmK8eGbS2ky1J18/Jvbw3jyjqtsAWTNime49HFirph/
6TvOJyZXGws0EPLjcG0NS8XfFzCleinB6uesBqsptGei+lki/ej1FgTEt1puD8Jw
X3WgpdMzI3UKC35aDhMU2Ni6ZjIcVaWVf4fdwJXGsu+heu0VcTWMnry3dABESMsd
CxBhPBTd8A9obQ7M3D2G4rZkXiGeCYfrQ2Pd99w8ZaA9eD0d/RayLLfwSd6pWyEp
RVfXCZ0Xnlfkazq/flzkA2pcKUlyEXsZaW6nM3LdL78pTV6VOM1sBiVj361tD07P
I5LOjM4KnzAL65iv6ax4FdqHxUoJe4hBeLxpm+r3gjmpyIXUWv31haAyq2yIaNir
AMDvUYdcnsv83JzE8QFhSa4IY5r/Pgi1P11oOL7tLKf7yurM2NWXEaXqJ99ueVqU
TdllsJsWIUNNI0wa+m4ohM9ZTpAqsS0bMk3aqHoV6yV4yiWdqbVJ08vXlADWVV/6
KD0v9FfPw93wyWsoIVSgu+DSFsrzjvbglalC9XKA2pG4l96TagVQ4pKrRyECNbEc
tkvaOu5xShBZ5j9snqDmY8YPG8qhcrGVyVQvmSigfgd2g/011YzJPXQeGyf4Z3Ar
SFvV8/rRKWz7HdZrFFOkRUAcITIiYD2h6VLUqTnhjJUJl/14ve/2LyO5IrrV2WV+
9AyTVqWrBiPhc+FlEzrOBC0h5Gz0Ok6mYYv2ka8LOZKouaHGNeABx5DBBJkj+Vdo
G2ip/odXGv7Qxqyi+9IPhb9FThQaakZUn3EksIHB+bbRDobJw0xXzltAb1PngnZS
mSL3Nms5YpcmHgxUC8Nbqu3NvQg5iMQt6JPPjOVFVHGsBpEDWeNJFEdKEmjF2Bnf
dL+DKvatnXM/XMsJvL5gs33+ahVpSdXvtv/Rq1MakbRjWWZLG7EqkVhYYqlK0Zrw
SP/bx0MfzXEkvgqJLl0954Sg2BWhjeQK9FRtwLasOlCn89TFzC85FMxziwm6fly3
QlEaS65hAWwPetZY7pD2hS5Zrxl+rysJd0EqLFv0m2Fagw6x7ds86NP5Q+T5Eo7m
uU18J2cTCIPIKGr7O/fUeOxgp7QycWl/JA4wupI3bDaBM71RP0Se+hsyYzz85cwE
A40hN0fbNiV/iiFtd+ckqM2uegDEklyGkXUrP7ZkUcq7WPfC8ixCjg04syxbIEDU
dQeHl5mySerJIlSIYzqAIEhseHeSFtdT18hOD1un8ra1Y4FMzaMzShMfpM0XxPFh
gdNBDkpP/jgQqusO9O/nzKmv78AV2/QcZwHabDY0IOMwY4uF74S3QEM71Wszc6y8
NFISr36oK+7HLoLIE6x5b2CV7UbO5Nvxqf4tlWPxavLJncdgGn0hENHCK5kOQTlC
aL0sXFnqdcYRYXulqTp8RLjIz2xkSz5d7qtmBJVajLjpuaTFrYLLHC1by7eIo6uv
HZOkcuzjzXJ0I30ON2IVGaWL/Xil5GYPeV+g1wF+EGMDqLQOOJ7nQ2nEFaaIox59
1JT2XI1t3lJ/1DyqHSLLrL41mVekFA/uxDzgq5GPhe2KZOGU0+39M05UkeX1pClp
2N937BeHL0DUVGfaw0O+Ggv+AVzlPf6kYFu4jxMQngSYW/O8glnlyae3XH73Pj2a
fXkW2PtXAjevySYfuDyfMBFDgmFsxlrGW5wLCU/Ax87LT7kjIkCLbOVcxbf/+gAx
wdF/FK3tktS/0V28VpKTNpc4B+tr8ldtiILo5MDj7/65RXzs5TrbHGdBUAbqMqnj
erad4rghjPbrDHOkJuVlM1yUsO1NsYV4nzit695JHKRAkdItgNUsWa63ZD/zeb7C
2owgC0QbkvS5YfQIFmTBeXOYUfUjrp1LM/rDPKUpgCMb/79LjdQ3InCY9jRRLyWb
fSgNt2cCmx67lSL7zmkBm08ja6OutjnudNrp66k4TZZrazXEqZcqoT00BV5gV0w7
t+VCESUA8hahNupHHMmotkSb4PeNE34b+UXpSvHAquioJydA4X7FMq15iicE0CoN
t8epCC1KBhBHCzbt3nwx1PHb3w6+8r5cBSiJImvPNz1+nnBScAdpO5/88M+IOET8
I5Y/H3wnGhjCVms17lz7UkLtk0xnMN8Q/U6XAYAR+UHtgMT87vC+g4fy6gtkvTIv
UDE+BKQpllLJyKU+VrN2TZOL1uum8MPu7DX+hEk8skBG6jlhon3c/G8k0zL/ZwAx
9PF8YJxcVv0z88cfKVcUsB8Uamlq8CleTQAUBhYU44rzwsIkvwkBxMpvikFLciyA
/+klG8IQePZuBIhv9hkdJGjg+sDDx4dCiuWhsng/VEDQQbBh8AUmay2BSomGbx63
CmygbAtz+O4+prJY5Qoe8GcIXDl6dnpqswoXcs65EM+r09aJ7hpsnU9MBwD5vBZx
tqcGRgz6uLSJdMNXJx4GGGt3+EdtQHdR7GvdAmVWKBTID9SspHztDL/akrNXjJF+
bUFl5Q0AUDWq7k3FsbxpHrTCFJehzPa119bV7W1IlSpLleMgwQcJocoI4fs3z2XO
i1WKgiZE1KVbyG/RERj0IuBbJmAM81uCYizTdoGUqPNB/lRQQtJNQCaTiOvERj7Q
A2bkTgFCZCarxXYF39/EHxXPl8Q7kgNcV1pHRY0Uxr06reUHW8UQ+BgbLeCUT1un
37QCsKrLHNzosZPkRcybsVXKFcuH+jHhW2fTYn8aVUnuC3VGGe0hgOC5hCv4bVVG
aiA5ASI0Bee6takHQs7rUpTNgyy+/ZYPnEyM7QWwOdls63YhZ7/a3iMxt+fvHRsm
thTcM4qFRMZDUb+Meww6NC0YVCqyFWBPECy0Zwax5QAkQgzSiJWJ8wWgKTv0jZjH
5Yq7iErbRPiA9OUa96AIXaQ0qGcwfdgJwdphVcS+o5/BUjYdEnR0eA0TFohs16dr
ILLW4YrKsuqUuqaGhqZ2pb6n0Xjj5KIfVapaXtAsPgPQHpZWo5ywrPToNVlPg7U1
+1wcBcoWLSAR7LzY5CSyNxf9QQwleKZyG5AUpuu7LodY5YqQ13xawLVi8Eag95/i
M2X4kblsUqF24LeSJTse45q+BzTU8G3Ecertl4Lb/kLKYGICBWAnI1GFY2DhNEoX
joSjNvF0u5gKEDhatsyuHgRYCr1/CKQUX4W2d0z9ZutWhTU8es1Tvr5GanA1L48F
7WSQdzcxatGsLiyQ0+dxDfmvxy6aatQXAzfHWm/nKOq1wwMS7rb5IRMUd4RTiB4I
fpI6pOs0c5RuJkLiZoCNSnEM72btWNM07ua3AEIEQpWBrCBdbTsoyaF94oOTkX6h
0jEgz2KdXXbOkt4b8oyEZ39LX3+NdjpcUVk/P00bs/lbsH70SSoOXklNyzWqdcE6
3y/olkRSGbA619S5wnWv4qqE5ijqKeGgIPXkumZk/qgbrGI+IlK9rUGFj36zb6BP
S8O6dZeoYrdi62IqLwDF8W7TWQTatwxnyfeQKXQL/4Zmy6SbuICsXjFJBhiOfUba
wOCxsjfBpgvvL9nRKnNZygUIcmGPOppI1D3tjDsMdEpRlbpP0XgQY5nUj1Ag2vOp
fxutovIj298ZIFrzqdxcIcrhe2RzvbeWpmyhEFNarrXan+oYYu5KiZJDwka4w58x
gW8TH9UYzG9vhHEykHObkyJLTm8r5MWz+7WJxf+3bZEwwwI7MMcS68L+nA7Xe2i/
lHgC/K/kJJ/vaRdnim6uyy84MmN2SWJeXmwFJup5+oxFH7YmKtUqFZEBbJQvx5Kk
xWHkFpvL4WZE/MhwgRA1QzT8jk4yiUbqvl1gc4ce2tP6JRumwfcLlKQPqEo6wDhc
v+Ah49y2wJIByh4LM+R6qAMacFa1gZZZqGL8ASk19o0m0vZFENgV7fK+ei6vfTS8
bwm2nrPjfarV+SKYy6e6j8/3IRXlZy4CvLKq4uZuANa/4eYlhP9raqoOmIkG1/Qn
B3flZcf7n+/fxh6tC/PA9it7WBVdDUm7vUbn1wxCssYXc7xuAe41QQz1U0wue7xe
DU+XG5wUKSmsIN/BQe87Wv5bi2JwMvUkhFM2pl/TV9QsURUud2z++zVm+UdQn0mZ
RFkqIgEq7PsZLSohNByV3CjMm8mJj+b+EKEv9FeQWNxLGJsd2RIn1nXJzb7qeazm
PPry5GbH9I41+BTuLVNn8S6dWNID7p++vfkUmkxgCBcxUPeFtPWaJlviMrGvdSdR
rA4/DA6cAob3SX2iIxMzd+QK9HYxb54nYcpphvTMKgdInh0yx4zbMk+k8QVZjs6F
C7iBn9M6DWlKw1gjLu7ZxdtvM7jINDeqoM7sGEGXFuA6JPQIwcx6NUeYIyKiAsBg
iH/S98Ti36Xkyq2em8GGcwrZp+rZ/ANPgE41C/1QNP+T6HNX8EnSn7mWL0EcsbNV
WUZu30u1VDk4pnAK1Nf9HsfIoDg8BamLMwuI+t7pR0XzPfAkmM05wa3X14ZdFxbp
O3ggh9AciuQyu0UhdsBXVtRdYyO0YaUh7SUeulaI9LgY9xkY+MGWkRrv+fDQAnP5
uexG2Vev3i1Qw8jhLXVYnyRqiyXnxL7nMVIZantcsRTsw1+e5wzAdMniJwNoKcNm
M1CmK3YB75W7GVHinU3kN/wNWHEt0UM9zK2iiKSCF3lnx/uFGWBtDZrLd39+GZVh
vFRuhvAO81jwNwfTC9titLqOMRZNPmaWpqsI455RuFTLHSCuTWrPPDdaKvoY64mQ
ilWI3PaGiDfNjcwSjiHYQEZOiUty/rqLPOII7gUMA+vKVDLTVhCcRNBlKbxzAT3k
hb91d9tM8PJ7/RC57Z8MEmq9MqVjlwSQdRHMyVLzkUbMENolf601Ykj9W6lVaHq/
Yu5+jFA0+kAB/t4HpiJFSC1q18PNS3vACenNcqHmFjO/ZNBvioMkjKTOBaTOzNQ0
oZHmSxMo7Q8XRQsl/Tgo6irus+PLifNrHdsqlzXaJA8lTf/t2mdOuOgIfpFtJHXL
o8l+PWiZDPmZbGJTVK7KxeZ4yV/XHCAGjNsPOyyo17/s4QjMdOCXZoJFxPDd1XCX
2Jk4Vg08sTnxTPt9830CDvLznIDpRgQY3jH/feFOxEt849baSquQiVS7K6yQzLsY
4niuLRpmpyycOQor9D8GTcBHoO/bMSnK2ugWC+JAOiK8tryoa9SI/XsSfZycCxpN
O8tzO9xT7Y/T5y2ryGChyWvyhPzl5IesTm3mU7/80tpiiNUwpsTFiKeoenjt0oSC
qkdJd2MbpxKiYBzI/WYrFJKdLVonclPL5Dfb3tcPI+gJYMXITlDFZXJyPKCeUUZL
x7VGPk2EnPzbKpWVyQ4N0nHfpTjqKy6yeB9tJdqQ2RmdRGajs5z1K3kl+bAO6E7U
X2lj+9h3umvLU64oGMMNK6haLaZC1rDQwegZtOT354njP7Xiv6Y3KYBCa3MYQnEg
W3ydPkXnaVELt921Py4oyshBQH/lmZEzB4lqPP4kyCpgz5HmqC7p5A8ry6CM1o8V
u81/wyDQ+VBDdQ8mL6OYUGhTbI7u1q5wgce/tUHKHrnOE/1YCjAkB+/mtgN1uy2Y
kzV2auC2wpc+bJjGun+hlwzey3EX4nFD2tVmfLEtlf2xCY4XDG6FmIz+2G5ZU9GM
JOrMwZBJGJ/y8v2CGUvE12BTafjKRZH8/9zEIEy6fN4yRBWiU+0sgQOdvmuzm+9v
XE2SD4BvC/deaUWQcA48j0L/dRxWnPafpwpynEpvfPgEwpK7ZWXdiD1TlMP2U+SR
Z0YO+g43dMj+44+UPwIqFLqjQi+DbE8enjbNpTOzcy9zpHjT0QkSad48wLjN2cIC
vJF/KVOq50hkJNpk1c4SkXjqaXUHGGQdsvPHKK5DAchqkrIR2615UJdk2lzSx3LB
BE6qkOHJ0Ct9uJSn1qE4XcVBJG3nSeP5ndUT+j57ej3WeXshZYOMqIIHLTbT7qFi
If0l+rRDWZHk5bQQpEPc2Ri62rLOXxlDLhOBIpRlN+gO+tnUlbHsRLM5V9tBI9kE
bDazlHToAX6YxsubhDPkooQsjmYpccSM6ONAJR11oZ3TTWwX84Q541uepLih69Zt
eMeujsreelZKDgj66W40OlibhQjAeouwZhVrGluvl6LYbjxYsNaF3JPbxRotdAZm
0E19b2vEOlwkOEwH7gvlSiqcDCAdpJLmyjN9HAtbknGbLo7VZktIWluFwNZ47Ytz
dpRBT4HlTwo6s8Lvi2w5cgqdgoLGBAI7M1umFt/TOAnWaxmBTbDDFCE77eyDY/H6
vECobBkDMFkdxqApKiRBroLXODegBbBAtd8L54JrxwITkB9NtaZGWXW8Kw8Kq517
Uw9+D9FCV3rCjrgszrRkdhHX0kVTSnBl3/0YB/1MbkbHhKv3JnptIigacxBmy9U3
hhuzfJF3WZ9XT6HKSHgQNHweFUmWRE+ECCiTyqCI65ftZrCOTq7UkGK4TeoNDOjy
vnpgjbwyYWvAEFskfCuSKbyRXmfYGfgKK3nsCSTugzc1tgQlkwPUAuTpwVCeEpra
Xfxxs+Fb9+g1IalCpRAvhbzRBgzqWQv6Ja+0GNmKsbCipvubnhsfcLHfv1/lW0LA
9Q6HTTwAwWfSkR5+fAKIvHo378qYBd8RAenX2BBjWHkEWbz7KDBBECNa7Q6Bn14U
tjIttLCcC7fuDm4YaxCGybX8iYdiYhP8WOX4IJ1U4ZqPm7qOox6W3EQUY3+2IAch
/S6M0zQ6rUJg7eD6St+migrraNoXuGZuv/fzK4+617CNtf8YHHP/VEcQKw9WvE0G
rbrPmJh/5TqlC0KCg5yhCAv7PRr4O6T7hyGtGfgavGXincaNA9g4z5JzcraLuTvi
eMEg43wdPZJOZIsJiGpcU5RSYlToG2Mr5IV7FtoWaCNlE3ibuGCfS5tsT1nAYUYk
2psh8oYlROX/HSIrleDNVlfF50PkYhnNC1blDrzL29NetiQTpQxmzL+O2GD/61zV
F1ZWeaanU3bd5KnkdxblRZ1wShElTrwHTa34EhKCuID4zV6cifj3SIwCIXE3xQs9
dSD116+HVzB4Hg90ZCdvD3l091E/LNRwXdTYjrJD7OErtw3pEjT36uXcuyfWkbN5
ZQJanOAI8BVB8k/DVIUvQ85LyWNCMgmHSU8k9qsUVt9Pdpov2X6Go1hmKpdY87yn
Giy7KDLeplzh7PCm4oMBkSu5WIuhhmwLF2amZNYrbn2DNkvTXKpRT47agV0a9/1Q
93yz87uhZF+mjID+Zq6vh71XLwCVDNOZHyWC0OkcJDZXnfzgSQbDpJHSIHTSwQ7R
zK/CYFyoSdPdgL4tfE0RqugZozgpxEHthIllYR9UVFzZtRD0FPfrtUcLhN73LiX2
sHjjeKuBMqK5FxAEU0TBOkyhN8LWWSAJJrxZQ766TCyaXL1VtFScVPmmv8Cc3v5Q
iEdEFlxHogvmIfVuyoskBldrXaGIwhUUtFzpefv3IXMfkdWjN2/OVMcRTshmILdq
83i598yO0RTZFv7o/EpOKK+L+chcGSsx77QXlH6gJZ4ARpztNXqaktict9DwSuaU
MRHeLPvu8gXsCgnfloGblH8SdZKgzxmVI5/9bCn4L39sVElmU/vVq0Kf75nPkf5y
Rafb1q8lZq6cx6w6JyBBrkHKC+2n+WP6UzZXP3MYDKMgO+gMl6TMJCCZFZHxpCgp
khu9FMfJ8gPVWgAkTtQvoXQ8MEyI64n9sdnYdXYyaqhKtLT0GL/UFch5hP1PIU+0
IFbW6bblvp/n655NdN3AeQ9l09K2kOXYQXpUsT6bceWAfFvdhFpyCVTbf/4GT1Md
pvzDbq2VVvzG7OAH3ncNsYfxBa8VvqL3zMxvxEnR9NULbpBogUYqpZcF4qDO59+B
V+RAnP/rrlfPdEGejmmomFSKPu+xhPEx4qpIdLvT42bgBiAUqzER+9joSLFq8ER1
JtfmHLG4O0qp9GZX741lz5vmUNMLFjugKlQqx5e9La7gApOLxmIuOMfXjjfpD03e
F2XJXNbHjNVdMQKpi1VYpbMj4kUt5ecVUzoEbDzkNY6fNs1KbXGkknQR76v9u0yi
zq6IvJ6cE7VFIW6SRr0Pu5NeVsx2zFBUO/I+JgWd6P+/eiXdiM6hrzsSeUqZaCj1
js0xRwj0fsXTHvvHwCb5HGLTo3HYe8ZLUyiRWTIZlw4TYQSaiRPUL+Rpnnn/l2D8
/Tx3TANEPB07L9HCBtdG3Q28eyWaGcAJgbyfQWRahWS83b4uk6YWGr9yVPDXkpLF
bie5dOh1QWizOUdzngq25mnv1LgF0fjMitH8KhEMrj8ldEm+6iwxJb8p+ke8J8Vf
aYIlC5pAXvmYzUtE1WurvELN6K4bzjGGC9iV02qe3jmTtAaV0SDs/JnoTpxbjeY2
bieOJ+z7AiGynntJ47yVNxKoks16BLSiqE84Y4xkKQngWBM1ga2umEblrGRzTtsu
QGp3U6hxTtLXyOpu66vZDaAGrV4MtiWXlsOEUiotujrdEWKZAGTkp3dSdWyag+bL
mJLvMPZ2JUnuoI1mZ4C8UO9w1mals/nhh51HhdyrzqtQe9Y+i474gfh2zsmibBkO
6xZaR/0YQZzIRpkM6j0v5WC87DzEMa6JI7mdoOWEKND5teEFhPDxoKUuGpDCSBYx
3lSI1b7xPhPKtLc/C1t81v6YEJD6b3A29WqtV2GQIpmZmuRhJalM0IJzSEESajPR
vgbH/6EMQYvSfYaJk6imHGpRc24OV/g4EI7PWcs4P7ljE7TBuAXuCByK/a26+d2a
67MNn/QmIXHp7zbW0KeizdbUHigbjYcDlGIeLFykndM8Z6D4luCu8uJLHT184WUR
m/ySfteezKEikXLSeX73s250mnDf/zOmd1aYegC3a7zlo0VXgfk1zivVeO+FrHCb
EORBQxhMSOS1pDgLJ2HKpWw7OFY62AaGJEjNoc28vvcIY6fDDVEzVfvcHIvCzqcF
Fr0RcmVz9uZH7Jmx/+WUUd64k5MawHl8UlH4DzTIHKVaiqZxRV20XRbga4xehkNZ
Vc30OareRgn0C8HzkB8P7dF5V9+c65FLS3uEgPeKYLJXIudDk4sFEtX5fpJ1jg/K
exZ3s1kM9fPzr14rWt9p7fj0WDziLA8fHgIcsyjTMkfVQy4poKtiKtV07A9PE49S
hFRpcEXajSZsUDtQEHl4hFQ2jWl5JxJwBaT2lihKUyTDJNroOvmMEYeTWWGBzxBP
iw6E1i8cEAa5exU2BfZTkPOsufgtrn2/4vYNCwGre2ZFXvp8hy8QBgdnD0m9D9EH
Sbf94OhuWUCTZr1cfk7yD5ltlz2SoXjZpTKGKQosiqAZ8M84DW55Hk/n0NcXzz7T
S17404CXwqTKhWetq6F/AtLhTlrwWeeyhuN1lzeAh338P+uFmKIJXpOh3edDE5hU
5pWhTAUlysoVLA5x+JhI6Y5HEutmYerjGPYa2Lur6KP9ndPq0XhogKdDg2/3OFxP
J/1CDgPZ0Ei28lxV8M+mhn+cKyOT0ySmdJqFOD0HRnCJnuAfm+EVNsU+Xjgcm+8d
Rsp6Trh2FGngYgzxAT7AQSbxnuFYIUTP2EMk6TDthMkJPBnbvn6XQlRHM/wmvYzI
hTNlyxQYpm6W1u2Zn6h/aztYVmAyb/y/3A8YcV4Mjx81cipmJ2wutM1+FN6cD9hN
UWI5t8RzB6ZhtJjhYfrZTrhSIL4FqXPRROLViFdMe39DSCd7rjldFnQV/5HOY2SM
lLHtNfMqRlnKajFFPK9wrCnzpmaFAdy+hsQ57AlY+Kze3BtH9R0osJ94IZok+45q
5r0PsrNBmQ2s/XhGAzkHwpYcEcbvYgq/MXOloKYXxiKYlPRNCu437tJquklnSd3b
C/9X+SzYJjpA8XPEBr4ASB9ja5t3uN+NdnEJ6wvaZy2UN1R74GpoKFv5EnDlzF2k
hU+x4miPYyxQXz9tx8yYreR7/u3Lry9esP74YmKCGfmA4h0Kcg4He039qifccxVw
LSz8tstX1bL5yoUsDcbjrZ/6ZHwar/PoO5i9bKkwcpuCMAKDnXMmnKKlMfYQDg6u
IJz1QICP5A+9yywBrTSoPNd9ooBNEgBYnTUbbgWGWkY/sYz19J2laGEbpD7Ypawl
Kgd9oCEAZsREDWJY5sgiFpN3/pRdSn3B4eXOyPrP3VvyFISusUrBLskDhMIj//A2
6+kGydAZTxGb0u0qvbsWxkwNy+y7M6DjF34CoxvoTTPGISBg4sHmv47F+naI8odB
FuZdL8uLZHVlxKcPv0Ka0zlGHBwpLvMPLPR/LqdVfT+P/O9AQs7giHyF9pUPHVA4
3CoEUrP7gRe4P/prb2uzI9/19lorHAvF+VYKqFiFRRVHnUG8e9+AQfhakuvcdZkv
QRsXuhE9k0aKaz0lHbH0kdMMF+rOQnyNd5nmdaJ4uoZu1v5s90V2noxFvoNagsl8
qtRKrVMF7rRAvt0UZIeEFh7pw2oQvVy8e9PGKV2M+CXIsebonl+5u2SBB0hZaVwb
6IRU0r6qN/WNoFJA3Wj4SEceA0z9sI3VXlTZbVSWdk6xsR0yZiVKKOupoJBboJWl
nuUIzHTaPz/7zGjwiG/RoXLHEJ0lKOohC+b49gWnHqOogiV+fhDWLbzkxiF5EJLr
wNwQPUiE4zftc6CU6s/FENi+pdi9bxgC6/g2FZaB5VB38ndbtYxM4KmKzCWxfmx0
KCTZW3SYdZNlZTqYyzjx6bPBwKd5NuFmtcZx6arq8Ix1HYa3sEVYDp/fGEnIj/bO
UWmkU5lCgPaSpKLR7DVas8Q5X4ahWmSdN7Fj4pKyTqzYkBDJv2bqtDweqIBXzv52
NJudTD/FtKsNOx0ueiESO9OfUtVpT0h8qs5vL5rHJgkYRKPYwx2SgUa/Z6m6n+4W
i4obccc7/XDQbyXemkzNAIzdV9KfOw9IIyPf4tsAMWTECaxdLChxMUFX+MlEFT7C
/FYUHwXStEX/LjmSpvqefX25nH6kmD3ThesGF4+WAmEiECeU59NJlzb+odE7e4K9
2wN+rV3w9QurQUavCvvVJWqS+8x1pO61hJ8oEd8WhFXbJzq//uDbFm++P4dRPA4r
ASdR/UNgMUOGP0J0HZetiOJ2/qMpHDj6RKpyT/+W7BDDtLPZWVvu/SLWgrDkTwUJ
1cGIS2sRE6YPlEF/vzwjkieRkbIVVp+jJNltTfjx+3yUwekME8XyJTnnub95KMTw
qDKh+I3gf6PNYm5Lc/WuOWVghRhFj/vVnXKVDLYY4OoS8qCS4zCNOZMYp7TNUkOW
zesa9myuPU1Momfh59oIMWY1S5oCxQF+1LL5QJRXC1j4tzRobJ+3UZPiZlaGD9Y0
BVPSNU4KQoj09aFhZbFPiwAOUPW5XCrQofWFfy6ZVIWtoFpstGTX88Lj+0LsBAa1
ANdLBNqwHhOae3LupC7LyW16TDq9Sl1z5H9bfO4Runn7PgOlspAWKkuC5TXnWVwj
FPsnlcnC89JR9DgdqJdmqCzpmSPuhGP0nKiXdln8Az9F34FGok2HAbMva4ya9+Yw
AJOCdoSKfOw8f7q2vU7okl8ka0IEUzqCTwI4S7YzGM1d+/WhSttpukfMFF3Tlxle
nKPVYn4XzwIMqC8HUT+h1TKgVl1dpiHzVpLeSUVDY4gLO3PVfZfg4Dq6Dk6Zky7f
QRKKsAjGZJEkqZpgaNodqXPhHby6R5lut0YuHDjEW5+0i5WknUHMTI8NF+hOsy6T
tZhlrLXJDKvoiWIJCXIzZRwugoyCIwQrz9+ZxSH+fnTQoJvf4QhHfHwbHCc6WPzr
qJtXunUG0RcZeNG/xrkDFLpTbmgcsSCv/pjAnqrq35aVQGbVLJ+t9kkNIm4Tpa+B
RgC5CWgUFViA0PeL9m9ZW1qej8FNYTGUbbWkNSX64sy4Isv2+6O9jMHf+jSKMdow
1Fnh7PfJGgTi44NwM6FAz6BZnnuYQp439AdKJa+KD0swVgVkfdBdXJ9Z/Xzr+AxM
L5Tc0Hm2cY4s7JimtVDpEproslsVG9sVEkV01UQT2v7HYvYVmZxrmvfwzuEihEGH
5aRhv1Yh+B8MbKKghYS5DNykn2F/IJkQ0x2y4n1aivOJ13nIlHYQNYFZZ6YGK3AE
XdVdc/HENixDAVnlG9jXTAuTe88z4dzb9dD48LBSc6hEjFBnh1mS0oeG6nnOs73/
LX6u+JxMfo5u0/IJuVrHAOeoTV5jErKtFTePesa+PkUOOa+G8Bu9F6kF9zZRfERT
nCcYa7FCm7AONRrzV4hZA/4IwP6z8hy+SWgNrn7g8eMXE9HnWR4uRp6WSazfshDT
K9AKAb0ueUvRj04pHh4ifDC6orZcrk2MRIHR6ZsC9sHrVLJnw5L2QmJLD7TLzQT4
7gPod6skTViPH3NDvX08Nq+vYugy3C4GCfw1u4VuRoJqdzcXJKLLVLcTvAKwUMTD
70tracrkxZIKfYfDl8YAFsSWN8U4nzGzgOx0TOJaPZtGu7AD+z2sCiYaLs6TWcB8
VGcGptr5Tf7WTGIMoSt7dPTKSkTHkVsNDS0WrTkS0hwDRTJK1W0LnhTFFFlROdqK
SX9YY2lC6J5BH6O/MKhfGiqYwXjcDCqURQ0XxIauzIpGib7aTigKljTrm5MLZw8u
FtWriUADfPSWR7UrNq+EpxvhZDPu3akT//B/iA4bQHh8g8R//f+KfDxNWHiaesZh
r70UqXfPhV7pVr1nwCJ9OovYEPffSpCCYaybIzhVysXNhYLe3ex3onp/6Dpp+Tuj
LZUFxDbgRu0k5OSUpvTkOYd338yq9LpTNMDCKYbd3f51zNLbfp1iFwZ/vTQ71t6Y
U9qK3pzN8Bt41/jfPtKBSKnrmuQ1cO7SOUsg2elxcqRtlb1rQVRIf2s5NkK28+jl
azL2o9YIfVVZciOwIgCmkSS8n6PX+j4TMCqwgOfIG+fV0zvq9o1yVUZPmbMXkuiA
rlLzF365poKZcL0qwMMg6slaaQFLqU3Nq7wk9HoqmH8QBDX1erFCvCTb07EP4Ib1
KpUZXqLzhkeH3+83TPO4PUGe+UzQW61TSubyX7thuMkZfA2b16OHrF2o4cg0xsIt
2zdd8Y5ZQQNnwcMT8WMVIzdCcy3H6bvVi56rc03siQCMN3b6BvndieG4LOQbM0V3
bzfxz7VPgc1czwonOdiRpZF/6/0QYwFhyhlFUas3oYXYNTHMpb+0QdmcuAGZDdbA
jhiqyvPkXfTf6aGMgvzixEk5krVXOAtFRc8V1H9Wm3X4+PXPBPAixIT8oR+cYNH5
/zUTVBWbK0/NEMYy24zV7ENgssXZukKDBk6xIVvb3FYgoYYY6HC/HtCDrakyQnax
ATfoQBMG7rqHNIWw0I7YcMXBdUhpQxm3ro4iqCHiDrj06MtTCYeSdC899myX6FuZ
z3mINOUg2p+5cAC4FgG7moOgv1K93u0C0SDuQbF5GzVTiTwpVGf70fMZ8N+nk/7b
3OeoK96QXmv+v61fXhdWWI74IS85z3uWCSFgHwlkMp6fiWJj9UK17WB0rsGb7Vv/
2DnUCnjkIl7dTcufOS+MXHM96z+Jna2Sphb940veOJXj1gwZgtfEPkPQ7ko4jBGD
l6NF6XeAlwxgcLq+gTj4/1rnGwQBw3tHUtjsKlB0QdASlbxDFebgxqXVFsDUJa9b
W+TDiYV8Lg2odeeMeY7jkzb3RO0akiviH1UEDyfjHIVkwi6IYmFj67/3Dt1ypPHB
p0CPN7V/DbosRWo6653MLHSQ67vxGdtGcl/Px8BqRf7H/ejGjJ9UpHLmZeVOBtjB
A8yE3+rf4BTkToHVx3GeSsY6v4ZmZx0wDK+Alt16n2LbFmu+k6c9s6OGa81Y07VM
eL+Xu60b9kXNlxw2dSA73pKkoSgXwlDx3L+vdfHpiU1bwiuNHZT8WF6dOIdTzNEg
pfFu+Mc3BGZVZR5FHZjnbKXXVdN+umhCCNJF0tLtND+K/8KSkndpf6IjoG9Qe2nv
DwDLni0Wu/u7KBzFbyF6waeADLe1RzQwrELMaOPq4AJbwvTgWJ7GI4x2Xh6MGHpk
IwYaedhhxeVLea0p3ZCmzloCDfG2KXoh8gDbADfBm1f2n2FnLQw4A1GiyQIvCVL+
yr8hU5v5/hTlTN6ujQ/TK5+SVyWv0eiH8Th0sd7PtAeKa5abJfsjh/iXSpIOsw8q
aALgbhLjNwXJZ2QRnmxAWLCAl0SVBv+BxcyTcSwFLdQWGUYr7u0cTRAC8KEeZ6T7
65c5Bb2vy4DXbg3s+PhOyzhOXh8kYpmXMsOcdCBkNg9JpWvb6fqcCXoESrLwBcll
S8qUuOPpAK4Ja5YAH8Cb5sBPjYciVf1fr+ZScywGVQaY/D6y9jwDPNgncGihm6MG
K04OvbGNhqqoWiXD3SWGadD8QpjDd4KSR9lxkKywMCw7Pytq7d71E/5ixNjPdHA0
t8NdZjX+r5ONaeKuzqnsopyyTkPBJS4/wmjWkn20/mnqBhLkPYxi9jVeExw5b0sy
v2DccYnUNOV5GN8BXmQZXzi8P/f6lSFF2Xn/gYELpD2Zpd6rt4B3V2aRcZVNB2vc
Jq4nd1k7inbjfRxpN75LVA5v62MgSaFPV/xwdlyhwmUZ9NfK9bvBKkm3Uhuh8TfU
YV9GcHJXUz0UXLDZe4MC9zUxk1hjnUquNBlKWt0wacSy8eozVY6oUa1HTGZqsORQ
8h6kf1pnAKeQqYEbTONY9w+694Zeh6HCrKXTM61XNlycMju1vu/6tSOgyMpMthhJ
S2b8AfJkXafmfqu2MKdEVfgSFk+L103iNPMHZNYlCfHpcb06rnskf9nu9KVQwhO7
F0z+eQYihS5wGTz4VOHieWnXfubxHZxVdxaZPLbH1Mt01u31AIzQZWM0/RXqcza9
8gm4ru07cfdpOBxncd4bqHOY91IOPIZk7LZPKV+uMyHTCCyBs2ZFGk9vbIeJhS1N
dNwq/+5aHlbcyKYsu6dfsV5NpKeTVHMecuN7jzerfBi9mptq3b1hBQZ1dgrZ2NE4
PogtUwT+tSvzwD8+0PbGwnAMu3+b4MvMF1+65Yi8xGq27ZnxSNtackqxDqHbqMo/
TjkYer2FViZFfDLUD6WkkWowt/1YEPGqxdHIWD+6QOWG9AXdZkldszsydEhqqML0
SVUcoY+zoIZSFxdnw43JZkswTGAnQx6BgFzU+MftFVcp3SwyuQDJ7QMUqc5/IDkl
jxYmmT9NFqhB45kAMtIMOrUNOAf6o9NjvXnhoGrxzYcEuluDfjxzpT6U41UdAucf
zOlJfwI9wfwSbS0ZcYJEqI0ML308BlOdSn2wjDu4/Yz7KlMKppN0KXJPdplNLLxD
jHJfk6X9aJQ5Rs2eAYhdYocFsAHl4MndS+dHgHDtNGevbFdH0ZrpafZYDuyTjtS3
OVJtmf+fYicoamxRFpof15Pa+soWwhmSloz2OfEYI5wcQHO01jADjEiTeLgweeI9
QwIc37APdt+QB3lNP9hQdZdaz1NBQKOU4vT8EKeNjr5NWAXNXkgb6E+R9J6Q3UMg
IB9y2VAacKfKtYHhMYErh8T7ddH9u+0jD2QQXGEzas6gbd+JktbV91eS1rwZ3FUV
vU5FoecXTJjGAVpDO52SkpqPCl7KQd3DqwpQi69+/Z7jATfyv+wwY4zXhJf8Zl0S
sfHmbPjK+HwTFr1/+LWrEedR5rv2ZfoV1OVnzEp9PHMO0ugQx7D86zx2zgFWuL3E
AyCrsoKfCbcHU+AulUdaEZzqCZrTr+aK0I/XgKiKmqA5ssOcA2CQufXkOPMobPfd
OgZKFnRKMBWH73jPb691lnzEX8g8WXKF6ms48+HCaCFEPlkVtG4oA/ftAhKEkIkm
YM+8G4H+LlJAPYWsj3OJserr8mnWSv2ulo+jd5rty1uTg6DDps4YmZOAIf7VuS5w
TF2erNRkEg7NlewDxDgVD7YRAJvPwYH3cU0EJOcW56FxkWY3Zhx0LTNXKdOHmxhr
2dDzJ4+52+4zWvJ82I8DHeNGVOcSnmqMyvPGhIy47n0gAsVPcLcqT65GSSkjV8TN
x+W7fIe64Ymwl/3yXQ4cKYPYaIAIrV+U4SbU3+NWAEox5FXu2d4hljAUkIvE5R9k
e8FILY3GIqRDzLXJVQTuwpeIqPyzFvxJQZS28Htea9Gcq4dUqGdeEhMQDWR/hXgx
JEi6qOInPl4XFeTGGo3O7fGRNTWiueHszQzdlzZGJhoQpvPOwA7lrjzsxG/dkWMv
WxAPGO0NLpJsWgOuMgNGETz40b+q7pJCHk+elbmg3+RfgJSu0YGKhVMo12e00bpC
FObe+74hXq12mxFHuPCdrxAoKsMNZ5dbG1K4iUTMaA7xIUrkX5BCNQz+NKgElZ0K
CNwWYUKMUQZheWiHUGu4yJQoo/UKEUW/USojw/MYKsH630imggJ4y6qjzDIlFXnV
7vkyQH/TImTz8VGfflhPY5gkOxWsgn7FjckkURGK5VSSmwJCFxD3s51pK+L/TEkD
Gof1J4mB10HA9K+KHjSBZfA6ySK5Lx3WtNo2NAt7V754wpOznvzSTBkO2kSV+EI3
3ujoz09BTRqO93nNVQ9tTQeUbvJsCVsCU4wgBWHOwctpsoQ5nOaMdGJ8mDtzC5e8
oazOJxeVBWwAs/yRSwNU/vK7TEmjy4yTa0Loc37erX0UsXFFzNOosKAMT2Gp4rbT
oEh0QNthXxZJt+84W3VRj1oPQQ42QgA//g7tfM5VmC++qgG5XvPEg7BbyLCcgQ45
14ms16fGZUhdiJ6XgC9NDzPltlyJBUaOQQ+GQ9GQMbcxChz1RwBBU67M23geWUXM
1jNscBHrptr6sz4mrfp5jtbbpZjAKGl+AvFAGacu3gkWmnbdKWZav6cUfz9PV7kg
lqWrpZAytVEAOUQZG0ITo1Of9K3O0rLswRpDgFg1WHEh4rLZRp9P2nG2hmLIM/NK
RBADKXOT/XNxzeLxCHE0ERSIOWL2NYB2EG2s5el5wXBuHfcJ0dYbB6MhKwRKqVnl
gSlWgq4uxn2rj8S6ycRn1pKFqCzNL69uz+1vOaIh0RdG/3Dq+xT+BmkwOb2+FWay
4BXGBr9UmiRZxCuP1bS72xcvt1qDY9kpI3745ppDmae7xvlI/LBAJKA75igPCCz3
p2lwOQI16HIIkA/L2PvvVb57Vu008NAvcg4RiB7dDyW47lHTdgSHMWkaLjoDvu9g
JYOeFMhHqXvrrA3B0vgCf1BPTnGOlnXaN1SM2g4aOTU7/1VzbjrwYtXvMBkadM1s
YwPLwo1Go2HFKxAQAsHdk+MeI1ITkpf45TmD1iGMypbFQzaoddQbbAdJ+toXkkcp
2b7m27B2Ff5pKVMc2ilI1tJ8GvwioTcsDZLveB3VYYpNfqu0fAj1NO1OpPAYbmq6
HfEH0QX/ctM/jrsy7+tFi1E7dM/Y0khwrnTd9Q8Rd5xnS65oxSocR1rUAIkt7FYI
p4yMKXg5d3Gm9NhuO8bfMVeTqWR4TOm8OukYatIcv4Y+st6qAMwXYhLNAKvWTD7l
/5hrTjNsEPyK1e8eGJ2ekDhF+a8XMDF9nLIMWV2M/FcjfBFsFmwhSqrUwp4jEtGF
yn0pwXMhg22FMP6baMfZzGAevy9gqcORQbb//pg6Tl1gQy/w22UwQSpJUOkriAJQ
PKepqjJo+U9tOP5ipHz8d1k/LTqQ+ReQhwXEo1CQeAqgs3PBtTeHHggJDJoI8070
tYYWoXqWArTJTIc2WTsxhlSVf+lTmxJpPd069mX80XzpTPamB70fZ/4esyUK9Ndm
GJ1D87D3UcDzKUAP6JH9XdvOTv4gJKb9/CxDOzTxeLCvpzAAd1M3+x4YX4L8OYF9
AiJpp0q4W1iYEqnS3ELhX2U5ik/83m56nN8PpfZDy76VjeNwf/I0hoGaps+pckhf
YtGlIR1+JKDuIs4PsYKJwKM0I49NFLh9QkgBflG3ss28/WLVkFKOHVBrI+BDLAye
OVFvIYhu3Hu9gXGqPyEXPZ6l1jvO6HDBlHWPYR3eixXsXUeXb81fGr7/NjpytaUE
dNtbf3Ul0sdqM/ny9NoQuHrczGkIacTRQdsOC9V+cHtoNqfiV5roviHEg6ObSX/E
VVm1cegkK40xxSuusMErXnkATOeCW/BCA6p2IDdf/7qKPcl57gIg9BE19TDF+01J
UH3r6rNsIwE37AfbYSEn3/c7yBhzON9j21JZvqa7Tl1xOJpWN00Njx7XENfs+dN4
qgy79706GJPSpQRpaBbPNXLT0wVH9L2jPdBCYbBqAoq8SbsJ61EnIrtMPKCzPkn6
ReVkYynCfeeQQG3Bfhl59Q2lFX9X1RF4JvkJfYk5si59Cw+6nhdO/fZKqqjB3nl1
YqNakfsnLfNENd0VOpyDOFGBpaxX5WJ9E3VmfM/ikbeCAVVPKSGy+5E1vE9JRqsa
YCE4sH1cyyDejDj8hUtEFeECr8ooZk5SD+D0Fb8IhxO5Cv7LxrQXNbBqvour3dhq
uizu7hLylm/KBScXY4PTv6bJgm/sBNX9pb4dRIEe0y7ECTgrmiRdFV/rGsyJhUMa
CeLjYP05WAhtg39iO7BirXekKWSt0AJKDmKTXo7pf7NU8mKVKzMKd8veNowjrgIU
i+hllvOhOmy3N/6idgTvAgaB+ZDg1Myb4uR8Fu/aNkJJnOyTMK8XzdiGFV50p3M6
lNeVTXR/wmaKri/CFkgxAt5oVz8ogJjQv2K78xQt55/7S6Ya/NsSqbGvMUjg5XlD
OIt6kvZUV5EHCzCv6fD0F0/W3EXqc2IZJ7DgqeMYTQYCS5g9AoO3LK/7zGAIsL6C
EtY/qeK+UhpZC9MoA66ZT0RxZl+iyI7VJSgdBrsKDl1TgUTjKYGSlPEkrcHDGwZQ
yYgaBlwwExk74bT3e5enqdq5KZtr5EQq/mqZv20wvLo6O+/Z5g7g3Zgld8wImzfB
Xn8yQcyQGnIahVek172EuCAJzpBQpPhtzXxmuMnc617tPjH8TuOkrqeFsQfLDpLg
fxn6WcXXxFDefwla4y4y3b3Bz6m9SnVMz4WSwxMlsl8+c7jn0mdzAY4v+yyPFvFl
0Xe4CDuxlwJ4rJGBERgtk3eRB41CigXai5KU7ZJry7fGk3tuAgl74tbkED9SWu10
b1a/n69GOgPR+sLgPRmvHX0FCNZhImaxuq9gMvsH+Cyxu9nIyWN8qxGtV4R0baRX
+2toKRPXMCbkl7tFlUUCX+wpWsyvhQOgnOA8bzfa0xSIgm77uvfW8Fki9Zjevy1r
SfW7l0pyXVHUG9WXqt3geS2mF7pzb/0t77tD6CCJw2XZIgAbsFqQZwrCxqQflkw0
+DCkb4PNy2THLW6z9DU9F/G5vwu3g6O5c0JNHKoR1nQoDY7xyeiW+EGjgBy0sU0U
GOEqNLuVQ75c+YggjtLwRprbx2Ga5E9hnvxkKwx+DtrceSgIpPYin3LHlVkT1BSK
BqWDVjNpdlEpqNK4on3i/XOyMYmlm/7UQjyUHY9pgX4swDe8bYSxg3qvi+Wmy0sV
Mg5zOgx8C70+cT1WqaT/9fXaNRslH8kZh1bubl73Eyn6F999k2/+DiUQCwIzRfxU
NWCpn1x2VlsTkQCvwWsvvVxMAMQUpb7oaCqvFR4Mr/zPuHuiwj/amX+e0B8zp+t0
nUGOnsYZlg3sjRHCcQnpvHiwb36DnrWLCyWRz2JlHlSvS3Y2Lnk3jj9XNrZnadAF
lbkY3syhia3B40yrevjAuPd13TUaWTCF+AqTZlnLc+do81RwCRgPHc+IHVnr0DGm
gwkvAhr2EB391A69eIF0SnnMXu2FweiFg2XMvMgBCItdJ++RZDo2fGRxtxJByPDV
TupRoALkeJUOewuJjYTDvQ2YG1LKp9vgkiqIMfAIsIe3x/hVkc5otNLhBO5wuCFB
fhJ8Xu6n9b7eigBY5H+kR+Jwtel9EPoAjorBGqR4tgLCgTkLo+WWptf9qV8PR1lD
q0BrjgY0/LNsTqgfqHTjAAGUuBziPu91hqhaCl7703nxUODFTQz/CgM3nw8BOxrO
Wml8v+aUWNFj0VBXKDiJLy0UqM7EnKhmEmnJFrA0or1SHA7Zlhs8I4k0CGxn0vEg
ROH/qRitr6P8xSZpa8L4EFZkEu9zebcB7in/6l1tDRabbngYvA8mD+hP6Otecxa5
1TGoGnqZudJksyWI0UGOB+qL8eEB9AHYZCmklP8iSnfee/M4ta9lVd9kXV3xNXyY
Cv/K5EDF/GVJa14R09hQ6+/Z5R3BCRHltcOMMrbbEVVkZpp3DAHwFYqa764B/tJV
kHJpG6/BMofSTsvvzG2Dlhc07nmGSBjRGwJIVbiAs4CgF3gvqpemOcU7l0j0t6MM
NK5U8Z6uwVkYlvX+LbaQr3zIqvRzMZeuczJ/TX2s8VCBAXx9TrYEPA6CI2ZveR5z
DYBClSHpz1qaFSme+uQtJrlMZe6eFGvo+EuCifowhDXWL6t4QIkif2ID4O32vCwV
DezAIFsIiQeeyUQy6ERv4dxi9Sg81Dd/SEIZaP06W5J6otFf/VxjquaQo6tMjzbG
9HRyZzu1kLpUC6iaUYyZc+zIGKjXDVDM9a0mu5k8GzMZZ88YWENLi7EkQucZ8P7s
5lj6kWBfqUUYujvHAgVJ0mdlSOX6fi5/QahDjU7ultk+BF6NEGZbOhLGmcN5lwkp
4D7wUwjFvnp3yHTw2+TC/43I0P8qHKcTkI1Hgu31aHp87yHYcXOOwlXi+ZmnsdHv
QdDvTEczAfI2k4dJYyDljFRsBHdO7IJNP2ZEGFiSHpz8+pX1uREtwAUaP8kvzNbd
YF/wYg2tJPZWVAiT59KV32YR+KVS+BJEqs3Pf0ZH2dDjsN6ufKoRdiyHDq8EXD4u
bsVptRTyZJ/WAFnndT05NGEOmAQpM6ltpcvkLekG2YLs8gguYcTpsJM8y2FbuvVZ
Tg5bA2pg73JzRy3O0UXjDG9uFovMxAbUhLFc+UVGJwrK6SFbmHEsni8Qov6OYWg7
DxTouH6IrpMaTZS48XoDguOFWMkUSAcibpOyb39BYBTzamKST89ePban37yOlhAf
7Iwji3LYfCf0nblYHO7S0m6eBDM8P6EvelSdSGh8LaonPF3+M30+RFQ+LnRkJHZl
iVX+1ILBmsHaDKRYygHZP0YvCc/X0ekrxAEsztW6FTu2o1BpAlUrwjUXJCAr/zsW
bkTCNO+7rfLiIh3NwgLgJBCBMcsCb5iBwhS9h7QsZGIjqW/mCsqy/sqSooOnRMDW
3V2cv1nu80S9vNs9azaY5NcgdbY6Zt30aTm467i0qpDHO608AgHXtSkG0qXgQYKh
oCaLEnnv8enHqE/JMvyWnZ2T47JSipcVFubAOZiFCdp6I+Y8mYU+iKi2J5FYyZkC
QZ+jmIRjQmq4SctPfObYxICf177EQm7x9EC+JK+6cFEOHyp3Dr6QJZaJEE7+jCvR
k2yFYIoMFZBB4JxiPaP+gn99jRC6t0+0tjYWg1W8mxacX2ZIBZ8OmEPLe6Glzy2K
PKzO2gaJtZ5ZsfbXAeNqZKNR4f8k0Tdx1SV6QQ/MCq9NNQhRTXq16O9Djf+BZRRv
CgE+pYInzDweZlq1aa4o1kt9d0nrl71uo2+xI9g51dIaPzBIesazfRCqbvDP+zFm
QhhVoMkCbOREznaQMYuVQ5oCqMWgb8Kf637tMWUPEm2UxE9NcuKlJFcMrYblrQXF
Mv9/Rux37q8DqFm4+WWfr5wTExP/1DMfApU1B83nRoKncCMCLfCsBFEnNOxqHMjM
snpsoQHHoTHYCq/JtFQtqnLtdWwcy7mG4lwR36TOLLwkPA/RQ6/6yjyNSQP4kKXr
N21HhlteAaLqJO3mThPNeG9zGLqvqrvVBOaAehx+29iDgNNqLa/EA0/WFyUFoIdy
ksWgU84FIHf5QpcMRfon3g3kiH5VjtW0wvdEXBheixUriKCdACSoMBEjlanae2Ee
YCUCyWLcw2yVGU0Yq3D4oAxMvcBzG6TWrJ40UzzGmJetmX9uU7hdZ3ZjtupzsedG
t+WPap+RcknVDgX+Jt4iyd1qH8XKO9jrzYjnhQ4k4zyjn3JOj6mtvitVJ5rhOXmJ
dKw6EvLZ1NgHfxdcTDsA34EZ1d3XwF96zQJgfPEbfC+yZ08kdcRH5AClDehThX0I
cItrA2MwCDcBmlZXqW2DLle0xeSt7Tsn1S/rcxVj7Ds4S5PY33TfUx6FpbBu+9Bz
VOtsC987BzxZ1EvqSWat5fjPjDKxzOMAuZ7e7bdun+6N1MpyWh8gKw8MI9oBWtnv
F4fYlcnUOjVyyJSpB0iNmS2zn7WP3hZwcaRtHx5ED8bMJ/HKLEOHoa3D//m0thQA
xNKhbbjEVsLMOO+v62fqbgmiJv6MqWSeWmqlEUnjYmhromTVahsG97IdjFxubqWY
5IlBqZtdJk7F/ujlLz+/29ggL9oGduuHmEm4nxrboqAx05CVsNgj3kYarLPfgsNM
QJQiC3LvukEdpUE28RLzJyV/TOm1GBlkCCuMLbgGibxp/jF9gsSACchb+UCdkih6
ZEmnvV2Zga4P2IboCKXNllqz+6MrPWDj4PX+16wlnj9HJurOcPkPtB4P0SDCs3vu
dFldT1fspLwMkeY/4FGr8ePubYlZ3vee2mudFdEfJ62RaneWySR7yfwbWQBoOuwD
1tv5xPh27ViFSHln3UqWPAyi3/6Zq4rwkWLpmOn/RYJHRqz86Sk3HgrGwZGcl4m3
RlPGeToocbwxJBEtFvFJ0aQNZkI4L6n3h82Te/nRMu2usahDMaoSUpxsSADyBy5P
uHGzKHrBlyFsbx1PhcMqC24C4Y30nqHtRpy7aVzdKtfC4vKu573+P1znWVSnem/R
7fT47Z/BOby4VRnwaauufSPGYWrAV8rgT/IYB3IcZqPKTs60A5vBHP7C4vkCxDaM
sVgHBCkYwu/S3qhdpC46F+vyS5RH0UzQNJnhPrOyaHbnq76iKEdDw5tZIt1eO5SB
aL/mfnmgTnQwrQ5Ig5Z2Z73/OW5+RKRrYHb34yhdDJovjTeLBkcZ7wnZiFw+1zHI
ucpuxni096I/xzYjbAa83MVeHVv4kACOzahonbiLYZxgHVGSXeBOunkR1/C0vdZX
PIPuqT3Qe2UQmI3aaRVgBp7aTm63USilu2wyPV2+GfadlGF70ACKVHaZGHwKNWVZ
wztG0coJ9sOXTQwCkoqmg6D+SQOUJXu344aj21+UR19bV/nhmDyX+15RqojXz90M
gBYzfxu20sSf6Dz6r68j479qsgjT3RHj/M4dMIf1sFtogCZyXVlWXAMVWjpHZxlu
wlBgFRj7dvrfXJ5ljjLC7ZOqlZrPZ6nECYlXK1McN/qlNW24bts+ZYqAZeAmDLHN
GoGy9n0F1MCYFw1BbThsQFJZx/EygwAwvIOniuYLRoMpqoi9hqYOERWYaKZB5n4y
VlAT8HHjSK+FeW8wuy1JmcpUl5HXpyC85VmNwa5vR0G3qMm8No4ZU/VoyyyosZz9
NOYWoW/pWYjMV6rJ6cEaWuHW1w3usJStnDHSpGl+PJWfwyuazX2qkTygXYqAWoiy
F8PuaMzb7DSJoX8X8IOO59bgjJ7nURUzXdKkswJSkPJ/JVsBQqt2DmGxfgMrS117
gc9T+VyFOMtWKPURzpI7YGzT/SMhMgW7AMRm3wAn8koqggDHa5ntI4l0qOQEKhUc
DepJNbqTMJHKB8AaHxEvtf+huBkSbpGArWrmD5Und4PcK61Gl6u0LHQSIIDm5bjg
mxsNj/JguMM8BksY18ACPLOOwJeKKVBsJ2FThST891+eUYukRut2WbTvMJbuNDzz
eh3K/3FGPxnUOh4Z8Kzm3T90aYbvm4NWGM/xCrgsK4+6MdPD7chUZR20nzPR0JV6
fj10pNxvwzmzZzjc7dTh8cS7WnG2gPoqeZH53xnXzSIkKK97ThM70U5BZ3O4wOc4
g8DsgM24ZS9wxutmPGesWkiDN5wchkgFTXMExfHUeQplr2zArxQ5D+zhQ83fAaO0
xCyKcTUS/7mf+BzXPNa/T/bQ3SBMX1IBpH1CqHgUBPKoLpv5as1IZl1uybX62m9C
On2kBZu3nFby6HSWo1QrZbvBSS3RSOrUFVZhVLS4ZEvXAK1eAgm+G0eyuWQxw1MQ
nKW7lVHDNgpKZntYC+Eqw5g5TRR3H09tYlp1tDPz6rdQJG2qAHqEah6DSnx0FDqT
IMYKXufAtoTxYkvAIVJVPXgS3bKCCQ20V40mcT5rkgybDjs2vOWSFCiFwoOR/Ffv
cSzj1Eog9tEH34SE7pqD9RcZVyMgi/jluvmzXmjoGqkxFD/D1Md+i/IAtOQ4wUzl
O/AFMEZeiyMpzmLs8A+sXMzK/b1zpKD9bhvH94SvP3iLMZ4F8q98ySaU0g9v64AS
cFJS8TJWxLsW/6WE7MhjCyW0UBKS5LPOhUk4UUOmCAAO9IN8vqn/nvcYPJ7W2ENd
ypdKiMR63L3zKci1eJvLxaIrwJ63tCL7HftrNioYKrye5yTE+oHfLd8wIm/gmcVI
G8EtVdsEa/jSSHopvmSNISkJHinas3TiNxhpf/dU/LJrmZsV9akyxs6h9Bv7DSOJ
t5zvZ3/doJDTu2Ym90yZmtDtdppKfPB2cL8VsaYVzQgy0oxfi6gGBjHIrPMbEGUv
kCbk1z1mqe0NRS/b5v/EN7ncw3SewuLYPHJ1NyF0ikdY836DtQMB9+J1U59WEEeE
/rIyCTvCFr6XG7Lp8eY2PVKR8MM5cqvMmzUXZFf1fRZR3JhJcMFebohI/NxG6831
yDFIU4VQ8CKuvX1AavRGRF2twg5Db5MKMJrzM5hsfsexF3LNi6ZHLrUUTG8rEe6k
nT/ffpOqV8p5RKWQd1P9Jt/FtJsYgE6WdbVNQXc4Dzt7+xEN9NqQ3o7UvBJQ0XT1
xir7y6PBm8jOwgP+i9FqzZEONMF34n2X/yVh5e7xyx2jMihcTx1X1bCxgIDo4hR7
SKJrADj5qY4Kwl4yUhZ69WF6y34+oN5cacMNMTG0YdvIe+LC3RdWDu3mMpgS3l7G
pmzjdu92JEfD9DXt8GMcj2i8ZuJb4yHM5viIW5PlpNtSVXBaBwC14TTd1UHuFums
7ZTwdhme0iqbweSC0S5oqrSMlKBkThiJfGtt42cbctZn2rO0IboRLL+RxUtZjALP
AASq2/V8S5PTeRwY+vWldcXdYMjPoth0b5BK5GeeNjjQTtZNqrvyMRbWPSQqjFZv
ytQD6/n1nPiShyYI1l4vPZplAwUXSmkxRQ6lI3aQ209iteGd5uwo7FzaGjvYKOXd
9axv8j5VJhMC4oQHlgUaE+HlxJ4nxvOiv9V6TlXsErAWnfpJAkAzelT3UCLXlUMV
agZMbUI7zHTdsIHVb5cXEj8IepQiLsoXWeyDlzuvrnuU8WKcT27ekuYK8uScfBTi
LOMb1XAoilnqo3uloNaLjeMZdW7fVaeLcrQYG5ljwHD7tq6hxJmAmhoJTJUS9iup
vZM1KoXI6Wg584vIZPOcks+JgxMiL2pOCTN36kMwlTJoELy3vrAQKfdiLSvgKYOr
93Od52PbEGg6G/4EaKWckDzn6MsVclC8GjfXn0EOvtj3L2mVeOC1e7TjGw9LPMjF
sGGCcsCHSlqh20DeP80euABPd7AePCuPfJlLntZmYfUeDnHskNZmbkF1TFZCYaCD
aHu8NdauBhtpFBqDs3u1iBVG+r1hXZEq69umboeYYdXKTJrdoa5m1H8Rbi+QkwIM
Td+NolkxwseRRsFASXuakh48EMuHS0JgxlIqLHAxG/4WEVmhNbIH7JYfSHABzATh
1ArvgXTrGpHK/IgF691RN8B2/qSpLYF3evhT0y+CIyDsi1oJr6MjjjvM2IasL+Bh
GifA0YNqihdlrvJ4Z5FZ1iPpmZYj2x1+QrHG1YpisnLfbsmV5DUdjxP8hrRddUwP
NL4tFVWCC1PMSHB6O2t07laNNpOikuexxr8p0ifOzaxjsqAYMteGJ20x0h4MiTSa
Xe9TeRb4AbUA7FC8ZDng6HTBdDLGRdC3ROJ63Tw8otFWXUoxUJKcwtYdftIcDuNf
IYO1mgIyjMRUtigcx0OEk6XB3XkPwNNTKU9M6b5BNNCndLMFkSz3AMOL380yzzKa
LZJtkv4W9+K9cOoCPbpxM17wOvb7ugfTepkF0/pj8ax3gFP7hE8ycR8xS43tlfth
KzncMJfFF5ZpMrBz49sYHedsaawIUHtaxEOeoS/SWOXInLrcPDW1V/SJOfO6biGP
wff34SdrE6Y+qQ0HeFIZZg+I1LhCuGfGHnDnHd6tR0fTd0ov/SH8bKNH+Qy/p3Kd
euhvbXMq4Kr8SCnKhs9yntIpiQqFc4EOfr3f/3vN2qZXuTZvXysj0vAI3vcPIkdE
apkNh0ZIQ233ICmRfkaRjGwDArb+UMsT7ALoM/OdCVWmPUGxHJUZTxsp90eKgnTq
/eqCeaN53lWhVBMZxOgsPg8s9KZhr9MRVbYpkCr/BhWLYM3qQdoVEXo7CALox8Sp
nhbRN53MbQl0uNz4UjMjRKwNI/JS3DOEpWBLOh+5jkEXDhjaV6jZNcBOhWRn7rq9
oncT/wLDlZHZpDGISfTCfN1OCbTNB+24JMpzFvVg98Gykr3m0hashcRNp7LXRTzM
a6fXsMsKCDAMwm/GNiU2YgTcmAyQSLCjqeaZB4qKU6PyVi6JpbvkaVva6VSIRS9v
LzojOuLaJ9Q+ItnW8gW9n3BIUntimWOMQ2KjriFUtOV5l5De8k4qljpxjfPjDaFO
0x5klEjtE2otu06kW6eeYGlqov5aI/5CNDuiCNKj5GpH5J1TYhmpdpIClo1YvdXK
kDxPk8/O+ZF1LstBRUmS+R9f1BPRLJPDttch8nMASzGL+Ob/VuJmo9xajLaD8CP4
Yo7MtZLcWAMx9USJi4W6Ryn74SLdXcsS0j/XacG4qFWiqnKspP8XIWe5qbz5d4Uu
d0+57LJP6u9hiVFQB7MlEXub7RKoSMiPhiVDseJHFSmQd+qCIe4FbUM2u6/31cOo
YsmRDN9ab42bbGBMrBBY7uBANsgoQNX4wWk0KYAD8ZzeJlydq+CqclsSZf+AEe1f
IhqxyQy+pNEQ4u2eGdD7sZDWFH1W/6ncUZcSQwrmsbxDCtnTJ4PGhk/ukHUr7JIM
ZE7qcQiM5yClSJ3YpPD3BTAlUmAYY2yUmK5+7vNTtE+KLlDEtUT82bycPatM22w6
B8XYixlrvgOjnW1QNjRN90j9KqXjRgkN2cbX4so9oZ2tdihmQjyIKCPlz2A/NaRW
BGjqcuW3rudKcvGX2veB03VRn4LOVuoSDoOaM7C6HZmXEfFvOi7Yd7OwHznbHgLR
YRDwPNzL4YRDA7ZLq9ubFTLDBLB4ARGN6BkRW5lockH83/SPXmC8uP0h6WgLBTSZ
E/akjaQc4NMMykX7HOBpJx19aShGMdBNpBRHZmkLo4kNQKK1DOEUaaqULW96/OZ6
t42f2hgKK4NH9i4AQ2BzLBu3OM/9mUe45+2MKwohQgWTKDzUQ+UVb7mShCDZTXQf
q6umREBlNL7JGkZvmGXO2iMMnKvTfZhtw3drsPtJA5sfrR06Tmqi1BU/4wwsYEO/
p93wZMWKcMBiK1ljj2XOXlAhnBFQbIfHlLOHuzIVMeRZ+rcvK85qy2BSPImpoGri
N6GVG/ZaMBlSkQTxdQG2VmfxYQ6Oa+G5Z8QmNSQvEd8+32VbWsH28D3FiKJ+DumQ
x4Q4BbCRVUrnnWCtuDWB7FOqGAqskNmyjKcAjxKx7eB/Obm7SS7tlQkZ6eBazxNQ
TV8dOWW5tr6BYmDohvh73QYnokK+zCNhlQDKv39kIGoJlSDJnnG7EOUgjYDW231q
MK4gJOl7FCLQlF/EK3xaNnrbN5RXsIXHeJJL9BECjUaC9suRA1pyLLehT54vcz6x
It4or8ghIEJAHoyLfr7m5LV/z30/bJhp2jHH//TS4z7JpnPGkblQHu0i6pHiYPaI
bjSCm2z11lQ1ocaek8d7+G3nty0haMJs0YJpXUvFKrOKkMnNSRfKjmUfKcBaVuBH
UulfBJ/SLAseMV6hOnXKhVi5imBD1OiQO1Vmbsa4bgQlHbF+5TV3oArVI5OuOaM+
2ZUKjHYzBWgv7Luz8dQQxhDLL9c3kns4p1dUl52NdAyAklJAdoeu7YOVRoeH+Ycz
GU2GY4PPQjAMKx7mbjYV1yg6SlZBXkayw6GtG986OsCSzJzLIErtnYymYCyteQ+E
t98+He5iB/VGIpkuMGscIQX8ehOhjcxs0WglP6sIadaoZfGQzFgmBvAIe5IVdgiL
nv5bfR8JQ5SPodI207bOlgVw0jrEFh4OWcbjX3iqf5wEx4BHXzil9K17+dQ9LVeE
0zhRQwuCADgAW1/JwYAC35sCYifrlr1ILvr7GjhVAWinjDollvK+/RvSou/Z/1XE
q3RkoDSy9i9RsKX2r38VLVtnZ6X5EDBiWVBRRQkJ+Ayd39qvnL7vUU2GyaxITUyE
VzW6uWo8KWumY681NjrZea5cRFe7fOjRIcVp1g6FQdpBJAmyQ31XWsBlamuAtI10
wOu0KyFF3IgMLRVbfIKiG0ptqrtSlll6wy5aBR3Ezmk4AGX8mJyQN0YWSfhbQDLi
DM+sud2y9slw+tJX7Qq4xFFtfiTUV6CbG4ILgrlX/Zdb3YJpS65I5t73zh24KxlL
hZMLYwPaqb7217chtAADlnC5IGg5QT3HoUYF6aEM+i8NtjGoB3uVguMAiC+/KY9n
mCaegecbA9ikrgMOJDDUY6MvPVoB/o6gOZObZV/lHsmvPzsbKx0tk1OsP/7r7yZO
SDGDRN73PETGn/7FkZUWvKn8yMe6IqotupuSKVPgE4ju3jUeyqelbnz9dE5Q9HFB
snU1d/4926GKPFIudjWrYlnghK4wXzeEbocBvzR8dbAfmgvr5oE1I9GOHNPoW2eV
GIuzKZUTlcBkGDzXFJRrFjqhRcPZh/5F9GNhz0ntDucuXDce8FjIaCSeVSfFxXOP
rpUj4azF7PzlCBBZ9IfgJORO8zDyGOZZ89AJnfQEF0GmDb9WDZTLEUyTZ1rOXtcV
bWblWWtF4LuH1lPcgi63SP8hqrh8TcRCVC7/bbsCrhYbhYtJt9h8812zh+EoS6v7
R+URuywRyEQoGK19Wc3IvNElHGqkCidNHls5fmQlIEUW6mJD37To5St+VBnIlZU5
USuaFHNg7bER8DYrn/f1K4V7121BXUfqTFVnn3Y7wQSaa3myIu/n6dVSqLF3da0s
+1rcAwqoqNCybLMUte/NVJIzc+9dgEYtENK8WEAjb7qcFL5+GkUUcJk1pOWnjr5I
1shqtc+NSxMeWY9+/4VHA+qQ+hNM7ofLs3IGgByg8EZ3aHUz1LgkxR7m5+dnphLF
A54Xh+p1jIiR5vMSCgw9XNoXireV4sCG0idOQGD6k+383n77hdmNS47iK5OdOdeu
wNJgRKea2XYcaQJ/ctXR/U3pJu8umdEpquocxAstHij1B5GbHkSj7INFScge/x+7
9FfnBhDLoLu9JsXT8Ji05FMstvQx+CshiDjBvKmyQSpKATTZQH+Y+10cwNwl1v9P
m9oFiTEetvyX+PLzAFPZh2hG6DSYRc2pyqKCAOKvpZsM2m2vMbH2VZCotL12VD8S
yuR6Y/ZpX2W4QxE3/T3vEUA6+I4p25lw9xAffoC2NQYz/vMBDDl3lT7hDAPoJ9ZC
vmEpSyr815EE73Vz6gUnMIpgm9DdbZ5f1iAvgeU2zgPjIipQEpTyXDzdMAm/r3Dx
bLDpqWSnQ0wpThej4GVOrGlIl6fLA8H/TDHyE7bfhonjqJexDavxrcV5g7m9Sj3/
ogUwV/YEL4BZzVywoBpIrS1NERcV1k1Gwz7IdHbF+JyCnhOgJy1EtSsXTBjP+HJ6
OeObKMvxc5QKeZuvOO1crunVCWwngMU91+s8Ep6rN/xrvp/haQmb5fFFp1+STVt8
DH/YCfK4LmVxEUD4/gtwc4qn3IoFfAIWHVHWD5jBji5biZx2XWsMfcB16aXVF90E
uwwJ5YWlZjoExwPE0NYNUMSI37nvg8evRmkx5Gp6Ox3Grv0GDH6c8CDQjNbX9Hd7
DqyB05BnVaBRLg4TGg1zsqzOiPOMp+ZbYv+jA17F9aH9Bl2VB8R4BM9O3ZLgNkLG
fMcNl9IwQwzUHxvnS8qnkybozdzD3igHYMet3X/zB8OfvfW+yH8SquA6B31iXDl6
0FnYAfqZLU7abf/s83HIIxAJWryUFg4ybWMTlY3JeoqfBDUMAJEoIpskzJP7L5Hp
LA1zIBxY9EnKNGJQDGZg5sxXveR9ovuxfJ0XKXVEHoelvqKX3OJlv6rj9UgZVtDG
N62TIsx0DQTVw4qsmzHgXCH2bYK/fVXKfL+0KmqjFOtvMKLAqa/XtmToD1LjhJFy
W4cS6vWD/B10H+hvMb4s+g5qzWKhJcDOeREF2M7iEgCcPJwam7UtjeRHJ9E5Jmhx
3hsDB+09NiWyzVM67lcc1CHaouiYnURPQpllUaT44LqgjpZwGzmUn6eTkHzwCZzb
+hIGD1n8E/6hbjzh76Q8JJoNkg1YRPGuZrtw5a/Noy1TZ6pCCkJczla1/+cUr1X0
MpEGa8lQpkqKhF9Bk0olDaBbBZ9RZy+GEu734nkK712JyEoi4LwuZpwMehQY5O+8
MMZxaKUDDuD+RkPAjIQetVt45d8som1qLVb+gmvrZMMy5/lXL0XwQGa+zHKPtfUP
5BCqWqYVOVhu2FEbh+/1y3yMi4oOmOqMJgTUemsPhMUG5KP5jmJbjRHSkyvgtQP7
m5SHUozA3H8CZRKrqyq9MHk8UjJdO61nPotf8YBFEn0KemG629GU31i4Pv4HvATN
ek791TSyBq05Tmi8xhSTnb0qyehXCglQPUnZ1AKspUb/C8Ce3gB5KP18+krKJ572
GtFaunI+uoqlDPpSHGg0EcLTYQcScUNdwqrxaonfWZZxUtrUNcEoneDGrdhXvk4m
Fma1uYpco4YUH6jDH95lGlhlOyVIkQqf55PjWY+jP0ZdnScAoggHAuEtr67H8oNy
YeB5t/cUekoVIx+Aky6VigPaZeVDnQIzl89Yts7Son99hjgP6p+H+2wWogxc1JjF
GHkE28ZFahFbX7z5CNwn5XmB5ZNcw2Tr0ZJojP4VdB2DU8EJbZrlTqDoACgUbGpd
tn3x3JROy08g+uZZpT+wcGqRqZuxD5mQqLEa4c8Ah5CQGHlj71jATpE0P6uYOS7/
EFKWmgOmxi8mPI0EbUdHhj6m+WA4irJE0M0Z9z8cPAPp5ZkxHAvPwQjpCvAFnHzi
6TTSNz+sMvOs+FQpBnvdyBvXG2JqRZPnHtbPavwN511IU5FUDtwVuDVPWBVBSUKf
K87ujoF+fhNOGE5RfzrXLLpWWhmm4jYCgH7saCnzJXH11Pbesso2It9xpExDnA4T
cIRFaBv67ec9A3uJ11H0wOVvbSaduMOETLqotULwo+dkNK9rZidgHeZl+9s945aC
CsUdDtG3soC/TzkPYCj1cJ0kVwImVyfkDhaijNWS/2VtXJIArUzaEwVVSqXbkY5C
SQlcNZ8JJKqcH/VjYzS+fWCkYInRDfVQyKONs+ke5IrnKIV1aP1RA39Zpc7tzPjA
9PcXizsxW8AvVbVwJJ06OsKO2yTB2LKqMXvy1jOLt7NVe5awCaJrhMGzET8WqhyM
SSNHv22APEESWX+ZMwmjpuznod8ofv0LaGWx2BwfkurCP9uLHUWueS5llMtLxC7G
Fj27WGxsmdIv3iv8wbHa6tyiyn3eJEt4Awv697o+JdwEwUcWL7MWKvwGVjAlTLoR
Byj5Idqwa0BhlLDRzN7vsHf0Bz7cMrQjg97t964AUnLttHokKHqUMFZkUcxaHnp0
EzilOWF2QK3R90ypj5+LWwnwpzR9ZMZRe3vD4co3K7Wwq+Pf6iK/sc4Cvg3GPoVF
P4XO7PmUBj/AGhIAXIxN9me72RAT/2HZMgXEUH601UeJCaD1SZ1Jgw5zWeRnjv+/
FylfPvLEmyVnO+dz6wwYwDmiZnSLHz8p18V75n+BnHXLHMkUuoauXGmImwr/3gFM
YMzl9YPabf8NvnO/CdIW0BeHxyfoRAlTJyJFHiz0p8RHrQJDS9sQWY0rYUXojYHA
kXYL5105zaRXRFVU0XoIF5g0CIMRvYVORnZZLK1VR1oJuqgUtm9p0Rnxn0qcXh7Z
AdeFlh/tzA12CzMzIOE1tsZz/dC1Xs8kondlyG+U9Lkz7fUskEl6O+V4fGOfVti0
1CUPrYiIg+T5ijtsCxUa5SwqDcgdo0I3ZWmpW4je1mg7Xmj1JhFZJcPb0WjqwamV
WHiBHakxuUey7DYmkPNAnQTDxisooZ1pVYjVguxLbD1BLw9D0DI+EWP9ocLnlqAJ
kwvSzsLJszkZvIcOypHIXcyTn3c3QOuPJk8J05MdQs1SQUtZ0sE06ctXFrLLu5yb
2RGMq3CYxHiKcz29A2/0OfaPAhMoS4PdJpFFV34rNWcBjBcao+ZMc+0pjJgsQbOM
fJxV3EL3Jyn4Wyk9RE3Qqs82oC3UxPRhhwYAGNpPDLDC+pK9zGfElLkVG9y0I79j
mdUSqUhDeGPCyBxN5d0RGW/cbgpEdVHmqJzdItEDXmX04c2mZp0SLo4LxbzNxR+S
73iOC8pHOuYaqLCbUWBOMOzh+/DPEAyfugvVDc6M3zA+lI6Z/+OzJpMbASqZmCBl
ZyikVDKhQq0v/QWJ3LmcYtzBH9FP/rDndJPTMzntr0sETuKSb4DrRkTetHLKHgfc
MY2iUcXJeHmaDlGEzem2tmfMVGyvZ/Jm1kguHG2qAYvm6EPjSslXbMWjTbVzTrEV
Er/e048pDVvD92aCv/CN2kIJJcGzNIOwslzFJWXZM5DeQ1WERjJsJuw78H7367Qh
uO5vtluhXjVXT9uoE2iOcvNwcur/CKRPKvxQ4uIrrm8EqegNip2/IZssM4Twy4dd
0AIUMF7R6DP1RCq5lfPDTvSaEs+2YsbDTguQljXjkyCw5ocUacessSZi/iD0qyfF
OfvVbls3/rYJWLlkwhpvtKU3qNLBoSLaxvLWAMP9oWu3mP3dgWpHPwPWYiHgU8EC
/db+bNQTA19CyAhJu7DQc5jxEe5EiohZgsSmspmr7vouXOKDP2Luu+w0CS0XBBpn
MT4MSjjrCXkFBUzGej3AQAlmF6ZNEixOBt3MwCRImrvsAsTKnf4WYNukjqtxJjcA
QioWYbGVlKUEV8bK68Dpn7mlPYOBXYvjTJfpYxu+c2+jZnZMO9clWndTHC3u4fq/
x2WKjPDQiyTDMFuVD5/nYe+7F799Qbce7pV0J3WFzdmhSa2fcn4HxWd7vc1xolil
C+zTLHyUZF0I6c38Y4qea16zG+Mky3d8hElXAqXYRtKCAyVeNhNj3bvSxrhxuCmx
jqm1roji2VJTdTS3XHIEIU9n9tMXFUdE8A9kzLqSTXOXdlazephVk29kQLKGw+wm
b8oz0vdIosCl6rvAk1FNeP9c58PgdgXlSCp0n/Z4tIgsuA1LZ1WVOsHH2/734wg/
y9s9KPdxGdm7NgpNAlrPqT8Fi7o4rfRIc4vpmyiuPctnlT/S6jHNuXsJEIt7ByC7
PDbCc+rIIHq4rFlwdI42Oy3YBsPLEiQELUWwUVgOMOiyOkUCFQrC464VwYtQJ30g
on4x9h3YBll58Wfu8dpVkN/qoKvtnmlyaK9uRvb+c1eydOjR+qhO/oybjGC9GJST
iC+EjFH91dsvsplx0Xp4GNm6bWGGsl7pJyIBdX+Y7B78nf1jFNEvehjbFZviPTZw
J06kaS35ylAfhBb/nzUsxUPYPR5oZAFkJS3kJz0R5e8NlfYBEVBm0C8Tnm2vloCc
B/OEp7jW60HpztbujludoNkWE0aoK9K+7m2suYC9oEUBwKq8F7QSnrU9vDaRgqNZ
w4gN067ZvTf2EdAI/ivYWFRb46CH1/iRctDpEgmX34po+yOkmUFSS3rzoDy+NnnA
vqqXnffkwGcXgy7zQR72WMCXtkQkx/jYPAO+PVqfuyv9iqkGxLpUkmMcmvOCmpCj
qVgDTIRz8JAhMzz3Ygeb3jnQkf7g4kvzvnh6WqmGdYvRTrbvRx1j9fT3NBreXSgB
c1O9h5oRU6MyOiUR5pfw4XiImIlOCOQ97OracgwbGTe2IAMVfxzt5yMFTrbZOs+B
clXBHDPk/P9QQTqZttFbFMUUowPNFKL8ztoe6xkvnPBkDolCaOuBEPNTPMF70+IV
i0YaeSk0uRjiq284JbXxOyBLyswxDxXNii7n47W6zDDjA92PvVZcYcT4hcc/tTJ/
S7897/ls6xOcjKBjVTBRxp3Kv5Yce119KOhxTUthTpuvdd4NH2Yz9aQAZ7vq6bPo
KP3PURqbJAaOnjIwguwcJz9ypdObcBdw3uEwJ58292jX74Dp9vSkeKlHOpqL+tgx
nIDUtcAPrJFugdrW9AQUW06DHtFyiHUdW4K5SiYO5HVDYpw3V1TX8OPBrZRfwvZ5
tpCt7+n3bBRQxS419ybMB0aCys1LN6ZJJRRH6oRxfoGlXMj7nbZNt52T2NLFd2BY
fvGGdY9ACRDhuYv3JyVWLhMOXXjT+L2g/hDaKePKUZkVHAbuh54t1G4jjvy29XvL
MUcwIOOGzW40wLNK8KyMu9NEK+gAWupTjYeCQdr1sf0kJ5glZ21DACpz6bMaGmKf
x8ATgnibRUgv62n3LhgfA1t5kW05ispxWiR/ivzq513opkAQMQQ/YSgCRhz3HuXC
ALnn0uwQalacNr+512x9k+cvh+3xZEM2feBMwMYmwrmfX+q7wnxi75WIrhH2h5P0
lYfRnwrVm1/bKzVjuCv7eb/RUIqznduI1mOsAHZspQ4wpJZq6yMs9iNs9vLkDdYJ
jz68ijbe6rC0YovNGnMqW1mtLng/KjD4h0EiTcTTXB+4TX2BJlFdut6pgp4KB+Jj
K69FnqjuvH27R3XGkxLqfsxH/hwgoE2K9EfOEQYYVdghHpop0psldIsHFuoeueDy
rN49Tw0KWrAub0N2pyd1+keB8y1/+3/hEVxiA2P6qttqPNp3YHRCt+9hUHv3l7Oa
MHAM/RMWGgaOf8B9UYseoRQwK60hhVZJRvCFEr7EwxfdNlKtmqCZBlFa5L8A9R8p
BsV1gWraQEZ+YdapW0qgnq00rT3H9S6zPBTdYfuWwdWWIYvMXJi8IVKMz1ZxtBF1
59VdmK6ROr0kwIBfXwydM6Yu2yQoAxWFQQMIvR45lAn6/YMNgb1tx1uGxRwZPI+M
GxZ4pqPW/rsIglKgDPsWSj8DdAoZ6FrOG2G7aki+aBsOYnzZG9XHrBI/zx/xaeCs
XdnYCd5BKYyXP2Fe/OlMh8ipocEAQVmlAZXnQrfyj2YHKPrNjOQ+xHTyMFJOwgrS
M4sIFM/lgy4XB2rhtLS5oqlmBe0xB6CGW+Rplzi8GROcjkQdtwI0KBoU1akvkeCs
S0YaHg9U3ZUb1WmcRC+wtuiEXNZi6osldiagi3dxRO+fl/Zn1g68IP8f/utEoFRK
bUQ0xg4poTycskDysr0j4xWF3inC169e2C5OHXCzPNP+Ra5QTfN5JsiDa27kvJ7y
XiSDcR+wh18boXveHbSWiEFG7K1UhsN9WtzDqKeaAqbGTAW9F1EAaZIzE7Q2SaSY
P51YVrMJSJ7qTEdonkyJSbYH1jZp3bhT9JkrqNTbFtBEKE0kAzfYtIUx0LaZozg1
6EbBS4Sme6psoItyR4nc1E8gZ4Df83NdeYIquj6ZVrqAyV/55NmxKE7fBD6RGH/x
4KSPPFCyoP/h+u3SwoNLGOrHB3bp+umY07W7+gbY6RB9ArGOOs+mmy+hJsLGojTC
zTqmryL3QjMvka0VOJKe1Xow04tGck+MTvKKIgvWNGa5s2N53lKJchLSBYrvvoUy
IHpkxRFL10dlDZ5x+6seWMkZINmugL/XM7rxHswqo6nF7eGg00VLDjjtEcUunXtu
OV+07ZSprkHl58+W7G4qESWsWFMPaXSLfo4K+fSTKgm2yzW3WWybTUbOb+W6jN5K
YE5Tn2SfRSii5XZqUAgYgeBpc9h9Shjy1HOWEvxGLp8C6DMv0Cku8CFRoI1Z1JOL
5tq/wN8VwBRIlu9DtTe5XBNuwYALEnGlyHDNM3ysqmy0cJgO0lWpmq3UCCtdXvEf
EkH+727dx2Uhho7VlV4P2Yqg2f9oAdD45K6jGYXG7j11BhRyc0bSHrRdjm79q6dx
M7u4Nxh3Y8D2Ddf9/zhoH4jCLgVe31yv7ZmYyIL0QXdSf+1XtrmTNZYBKx5HZ/8w
Ny6sr5csYSD8OqrhcKWCmkukuiZQctUxfur8BjjC4coBht/GFLmGqTOldoTfTlg7
Y1QRkQNKEqJO/ZH0PRw02Xe44fZDppIyyZA3pyqPZtdXKdoFqVULruUvQhtdYoDy
xZESohkEF5/0ux+T3AFVKRocaTXs5WFHhedOC2QwWfN45kLTG58E0yHUf5H301+s
3/wWIzUYtbkjxDbBjV/Nd+2pQoGf7/29jagX2pjegkuACYhoPE8hQ8Qb+EeiBAYp
+moRgdVgO+98pRDyR79wZ/wnQodGQFGUKDwZmNaGKUJkyAc+qN+QlXZ+O3Bni6Rw
hRRVYdxPbeYFZrO11pYtECESNhzZXK6hmRq62YVOSGtlPJX/D4++5RisyD4Pu2hX
AsvkWNsP6s5CQGB8H6oxPNgzOvBWb8e6MjG5oU3C/UDukJlKhglbENCsuF0zjuJT
b+5BpZmEx0WLnHBYvbbyUwcpJ2O1AiI0tX7o8NEvcvDIV7uMZ27aqeLcVVkLdWis
GJro7GwWWDRfBbt4evdTLWiqGuSBUBVSW7bjJAkKsNWD+axLZJI5/C9DtNCBG+bl
Rcpc+7MgpVRw2dOXKFp7VYL0ojFYyvT2jUqx0F30qs8fiH4ZexleAXzrPARmkyVG
uMqPLrGJukL0Tn4EABc4XRU+rzTOrvoKzKNpNW2n/3ntWHLIfJoZsCt5AseoEzsJ
EHNpoq9U2B/pEAMS1OawkXNvoKlmFTNwp5qGmlLoYrMTf7+fdYv9QwsWOXTL2XHh
D2novPzaSxIqCSuJmmTLFe/FUSNB8DrEvsvrRGWzGfNRBznJStiKpgugiaFcExF+
uEZMsRExAwU0oFgL6uwUWXM5zFA1O1smPwtjl+f0WthjBrwVY+wN2KpsotjjkC/y
P4ZQ2Vd//jhZelI8BE3xF/QLDxdB/FpskzCaHVOOfaEljkXElRgxUy4iuAxsdiMH
AnlQ9ql/OSzvknZKR1WQZlFP5vk2F+BBgdT4jQvGk7UI6owUQqC52quaNPcBNdWz
NB73iDfg4F04Xdz90LQ3H4uGk/BPWQK77nemvM5Kl+RdkBZ+Hbwb1ri82ZXnSgHY
rBL+SPus+CU+MH8lIN+zfh15BA6nEPwQrMU2peKK4YVdihw+c8nmhqTykKbEcS7i
aez7+O64xXsR3WPKmx8MZl4h5pTztKwksBLzIIc8n4CmbJc8EuC++csU/EjuSQHi
3XxpvWYkDBpCR8XzN50IMzx++Ue8U6aP2E7SnzUhhvDR5/OQfaKExJP7LAOAYzyp
nCq48772uE3+6QmNs04f7KtiLhRJa8ye2r8M+qg4KZKzuorOGo+XDJ1+h6/vQlL4
ZEeuqaKw/mhXZQfkgs0pEsH5iI2AUVut/o6Qlq2X/Ee6/IqNG2V66r3ZxCli0tDw
Il1+Nzaqnwka2YBbb54pqCQRhVJyIy/CNUwa5Ck1sQUgyS71dcd0ieUiA7hG7PLB
Jr3lSafpQ9/9BE+4bHcwILKNxffibP8RIUYze3uMWNKi4O/vwS7FGOdWBAjaVfXT
1gB5JYMWC6YWJ8avSLWZGIFeHYbXReNl3upS0ITRZa3NDJXYD0U20APPe8nPX/TR
QBlrcnxoc0SXJ+nQvIvCFWLI7uipsnj1XO3NNW5if8sIW3Uvr7y/7ct+Zeyxm2jy
HhGANI6sMJt9tjvKA3CGgokZt0+bfw71Yq4eOsAyyi6Bhds2MBC1D6uQFXg4fCbK
NBRAPw6BhMSIiOcaRIqZj72EUJxG+/4UCDf9yNwmXusinUHgOT7Ie5vb/P0XxQOV
CDZz8vfXYnCpbWB5qqdnYdbxYfeFVUxcVHhcZTz3EJWRgO+O/3+IsTBR0NXxPES7
tr1ElXBm+qlw+nCh9u0j6ND6IitSPjn3/v79E6ctOCmOVZy52xUI6wrdsO/NvSfq
/y81OBioNTTCNw912UK9RIwOELJQlES0w8BeyRnUVIhxBX5dfY8vOayNPvH44lng
4y6VsEuLJRPvC7ptK1EPNneqEY/aCTDjJpFvu2ncFSVUjLgNH0/KLLrV117Q6zyv
39a2WRKFDfQqdfkmH9P7NL1DgdhrM14alI0PQUYAlWvBc96gNYnQXqEgNmHGW9x7
07hE40g+o/X2TM51zNvVBwiIvqDshetIUKMsrMeS1SR99HOTP95OPkfK8KtjwzxN
pCQYI2HcCvsOyh93NzqEznQyj8Xa4jAlNcnz1lanAmvZ1EoMMjI85WVuz5kgC6d/
Zlg5VxgBLcS4DjqPv1F6V0GCSyuWtPwGBEj226ayiAkYidLNcMIZoG30PNc9YbXZ
o8dYZCOwWele9L45Y9voiteOm6fkM4lqGs+PRj/gQVrPb5lIn1isZdJPgE91WDyL
9QrNssqy5hYenurDUcbYCVSegQuXoEAbDHvaQ2wiwk/rmY2tNOY6pIzyGOIwBoCx
0xJ1pXWKQQULymQnUsUk52VmjWyuNe5NUqHCMjShq3VPljYCmzJwV8W3qp7P6LPm
8xOBh2baWhQUqlUIKGzrGzXMgc9h6mmjVh27Of54L351oKYbLLB/SAS0ZHPQGD9J
OF2wAZYgqpdG5np6zLCZ8gfbMFKIE6CSoOn5kgDfQunUO0fGDVbrqSFz1KyViIbP
X6e8NMSuCT49VA2gATNDtISkEpY3yKqvbYKZvd5BDbo4GhuTKX/+jbR7+pMQC41U
SaTJjQ2rkibx8B9BiMOe2yM/JHqQ/ql+DumpQcLtwWb1TeOtL0vUd6yIXbmrnjGy
Q7IBmPvDee3dwUnXUY0dOaMJ4Ddse6T1+2p2dZlgoqRgfoGodzr82W+tr/XGpHhb
KGCUvmGSkCOjkimWk0bqQHeXZq53Q2KJvDE0hEC5WQuvVD8/N2SuX9RthJI7KjGe
5euuToaVDIiY6XvelzDULDceqyWBhn8EaEnC7AFXOwPgmuNXELY5cjTdDSW2PVKB
9O3h5wRHD8CtWNqKN1PIBqA5R62okheEKPXDYgXqAlMby+eUDfYpGGcJCRoDYtYi
eI1Y0ohTcsVh+XiyC2WBBKSsOmNNBp22bRdmT9hK9ejjdg3KwXccy8WD68hKNZc/
2uvCDUBy7yXt1gaf6SLak9626BmzQv0+lD2Jw8wS4oavaMThdGaNeZhRHuy1TGFa
JuhfAT4UjAsRhA1pF9JrofdkJbOXyLEhpj2AJsUcXbbW5wWr7X2TlbduKcYEmrKm
bBchtHYnTXwLWUSsNIyGREWEue/va3e6AjW4NgFaCYh/YHRYuEkq3Qs5+5P7/Jsb
L5EB0Ar9Z96wRAQwYRWtKDavwX/g8fLqJ2cUP3hHEkWDQ9J4x8JpcREI2K5z9ctB
3EKYyASPFM6IYV47M4Z/ILmj50Ht+Wc6f8X8LrO0p7LvRAlLvUDZj7oTjw+hqa/M
+UJLWOgzY6sUVk94DcuxT7v18mxqUm6se2FM/w8BeLSQdzhdgEy3oDniruEvXEJj
8bGtp5fTe76UoMtivmgdTfaELov1yJ8AlffbBj+7EWfK06uxdjnldMjw2Kiogdgp
/TrWWl3e+2ANU7OUJu1iE7PxTTbRZWtJOb/AmfRXOLI0DrxN5Ob4mccZN2Gqc17f
/KbpnVH/w7XMeB40dQXgzpE6Wk8Vu1eZR0Akgqk1wcz2I8djLPWxgT6EcRps1CHa
BFka0WHjkCjSVg24caX1J2ou7tm0/XuhDc+E2GDmJMIJFB6dbGi3ubRyCldddNwM
YWHTeOCbHaXTcB0ENNx6/rdl0oWbfnoICjYizTI1dhvcO5nV+ZHzj/DeQXKNv/Q9
jUlPeCIRhlmLLwvAajnRHB6oresbesEXvOLRYYlZLkVuu3C0Y/CbUoacrAXhiaGa
NFi8DVM3UFM6s4zi/mpgfiNg+QqmCfkSFiKFmcguRluhhS3yjuEludrl0qKpA9jz
zfEHcghxH0wdFOrBT88c1nzvFjQdnvA/whUSvhejZRjQ4E0VMBN4Zf/YkNY21zBS
tWdBEncr3fytEHUI9hhu6fh7zs67q+34XQL3JGgdKS8n6/4PEZMNUgvLfE026qs0
SKfSeG6X/DHk3NY3te/BS+0VFtuKKy1NIrg2l7sW2N5BoondYyhHNTeBS+xcbtQb
LfODKToqpsKmsVai8wS8ifKRaR462p9GkEIoBNRzoIvbgFaEbxgnCzww8rnkK11+
xcfs0UfpL7w2wCcRpBL91hXtPrbcqNJTdWi3QFBQh7E9Bx8Ls/j0Y5s1SuTWcnIV
SEXqps2H+67Mj3NThQi9gyxYxof6gXS2yJccloNWMPr17efrl2l6V3X3EgLO0nln
6BL79cpw9qlOkn76CEmFXcMtSzOXMQjq0zsYlguRYIZMnwsE8ndP18oK8PU/NcS4
0O/yBA7mfTTq6KgWtFV+m/IF1NUr7lId5qBZqYLGisnU3gi03ico5Uz3J0ws+pgn
xlobTNmZI1HIxO114wWb/pjirEREIJoHNgkxaWP6lG2H1jS8NgfqdNZL+4oOLUbl
VQUPIC58ZE3cs3VJNwAxskMqpR8gQ2rTHdhQTdSHDuTdNCPraTra9/ozBNZgx7KD
TVrOUiMmECDW2B4MXMeBnAgyyDenwDFtuF9NnF56b6G4/NPcfWQiuTtCAb9i1Eby
F+AhOW9oV7qkBHgJlWwxaDmy2ZHw/ePDxicb4nhFhYCpXxi1e+q/RJwJOvXfMRcY
0OM/VuVQO3j5puJAKsfbOPYXgKmZI/ud3CdG/yAIGpDzWXrafbOJyVaLnzCsC/uc
+MeajAehGyDnoMiu2I8PgY5dqr8gZO29D/F6sXrqYSHuCNAFlopVlclHOjOcb6wN
BHh2yQeIvWZ5uwVNwtW2SIEUUeL5lniwRU33KJVtcUW1EAcJlQEJqK3Cq3lUfmOT
TgSrybv/O7+QzAFkf5BmE6gtQiEzjrXYCyVTRzkazmULmvHSAZy6MfbMYie0bfao
4fq9aaKKOo+maWtQIM/IGmsb4lLL3uFPmtZQPbnioTpcAsoHpZC+L1HvV2RkzB4m
zxb+Rxs2W9CS9p4aYV/3Bm2RXunG+yL+7KZHteeTQZoo4DzNOUQ2ZsqGgpzk1GbJ
JVlQgvuODnoLctGtdXp4nGTQqhLoI30ZBn5gOfLbcQumJel5xir7SXA0zHH04qo4
B1jeAtrbcVgBmnzCV611riYQ05pXc7sMjHwxrFMK5t3xzdQZuOR44Iy/3r4s+c9D
lEkqGpW1wVqgvailCUHWbipxbYXt1MpW1q78nCfaPm9xPz0upviPwC7jO3WzqY/K
M0VnPlZEU1g37pNglPYqHjnTeCoRzOAFNFDpZ0ZyI43C2WzICxT0grqlslS+ZZwK
3WchWX5L2/itv4bjN2Dd00w4oCYBjLynOC18rRn++Uir9MZ7SnnxW+8sCV3mEa80
0g8u+5qAvpahshGQqfzyZCwqX6g9a7k0TdCQbHw4VoZDSSN5np+82HNG5PfwXqMX
P32HdRqxmIhxEKnPes4PYtdZrCdSxV126lbzmayytLjM7FELtEvhbFdG+wohMTg8
g037d9Q6ZSiVcLvH2jBb9i6Nm3yK0qIEIZaBLzEldpnL91t/4J7jeOJ1UcP07hfK
Eoonxryz4GIJ4b8ojbUWghv5x2Eu7Le7n9EAckUmRwYPKcvjjl/Sqw7KR1yj653F
bFBpbX4aFpTR4nMMWa2NNV5uCyoycHmpepVfgKx2W8sSslRDC3UTpEEa9Hq9VuF2
DGTEYgS49tXZ4RaS25IzmcS1Vk3H7PRKphow5UVsteSJN8XlF8bb+q4GR4voBf+X
/EJaI1KQ5+ubn+4nYv7GxPCfpn/ruDCzK2jvP449OhXlDr+Kig0ZPzkUG2tuMnsR
mQhmS1GKqFPUls0lRvmax/ul2viM4IUtzx5lQUd/6u8YaZlzlpAntbFQmxPBM1Ha
046zLC2sbNY+FR51qbMC4GY1rHiPuPkxlktk4Tou+OBm32VnZkwCbsf6wG3Pikq9
/IGnNPIBSTfyknLs7wfMYD917ku/kMDvvuGKFfHR+uY0YADSMHwd7qHSzNcQ6JVE
2ZrgMCH1OmA6MfTJcc9pLnyGleHSsz5LFGZ8bN7va/2smd1hkoTICaV14QE5cABr
SIrBlOUrPGOnAOhNm2DyPfIVwrgebzVuXgHZ4r4z/LpIA9jyFWclr++pFkylxPTK
7Ndu0kcx9OAbrelBxdxSmuXI3EjNLxPh+j16goDIHN9kdPstWMywvYYILGbw8od+
iuF74tMYKMfk8B4xUR9/itur8CC/jFsjgdMvWsKjpYh+9unX7ayPcqbRr8w0h7ID
xSVWnx4xGYVJTdytTeUNnCorMA2PSceWTArMtIuoHnwpiluGz+R29qgjuMSlbh5s
WwrnfSyPMG2e8COu+SEESSjMZDj2Y5d804nSAREUTvYy8eAl5CMpvY/LpEGzduf3
5qxMPjDtxZs8fLvsfMcz3KjWO4etHgzyE3FMMDubTeiRgqj3gmKN8zEhyeUE3hr8
g1XLCUVBtWDki9YQUMJOk+xR0T6gUE8+3Xp5mVowTdP3bxQ8LlWjXutiMzU9fa76
imgtVGnWOWsrdh7v5NI0+A4IaKrp7t7u+c5ZOhNt5/vYrds9vOAyfPSzWnBILYV9
Y519llVyh3qB+aCL0JrTowLXOMlso6o9clxI2VN5z53OazjT8vpze9cATCAc2cX8
EInG2NoDx4TRiw3Jw0S7ze4mVXu6LGCBI/67SfzllXiGtD3UqWiAfZosjLMmesy2
WxCXNpdDAQYs8TvgaNQr4C4oJA8Bc0et/k54SJwj+D1PehgWbgMG7ngGu4ksPrho
FtxpmeMq34uRQ5p1qBgbs19zoCqXK6ooM62m1v3ywmzOqOHEx5uyqaZJgdUuPdGF
s5TqOGqagnVio9wKzFHuSrzkUneC62bP+heDtq5bov3CrDmIyhx16fio6V2VczPD
JVgLLlWVdEzEOaNJgNSRM6GhuFbdWqJK4jkhwaQa8mk/+YWAdGhlDl/TbWSSYBis
aPN1gz6WlaGrq3oawF39hudlue+rlBWjv+tSFnDbJF3Sg7xix4FY7UEwBCKbRl17
010kYLAwO3Kv3GxEUiePu/OEcCjXFw5z8UFmgshDSv2tw5bCU7d7SEJnPLO0iYWg
BZSfmQ1rcqlIZrYY/6ZtkNEIn+PCCBSiaTvQairvDWpwtm8wNBt7yLYZeYXlN9q2
6w2CTeZf0qiZqtD7Xyyr2WMq9T7VL+Mr/rsu6sq16y18bAECCbQC1lIGoJizIzpC
/vCa7sZWEF/Qr/LN5IvZC1g32829nYPVuboyn6F8o4+LzngYCU15YvtTvMcmt73t
rZzSppduUKIYHjQz0cdLeQxgMuqhj3MlJXkSRlJNgBe+39wRLOi0WjWr2tuerhnw
Bab22V6Sww/2lZJgj6IiwqRqbAsNi1VNkgDtp8Et+9lvUjmcrqBbbT8E+3URsG8n
U0M1Cgy5DgYXoaS8KaDARNviMvSscDRq8f5KXLEyAAS79kyGzIbn6vJryJJi4DkO
mWKmU4wn5Chn9LSQ271ITA0JDmNCPa2bQmMOCKt81Yt6U5wE1EqbcLsfEaHE22XZ
+HwU0JzmrGsz2VJNYA+ufzk+g13ft0+lCDW5rt1i58JmQRW1YfX4XnprF3urQEYZ
H116QZr1EJ9j5KAY7wj9RESshCIcNtkhxYi9TjG/Le/lXlR8R6gMk/TJw/nZpzUW
SBdAof7xvRoPaJNudlZEwJzMhOVkVuwMh3Xm9zngzO9gcREuaYNFVn33TY/1p9l3
rKoRBKrODTIcG5vKH7Tr58oxnjaKFXR277SRbLmsGzmVcHdp6rh1Eqxcz0qGS5PU
tQjJ+WdnFyQZTaa1iMd1gnb1E9hfURXy57isfSUQd/vElv73jf9yDzj2gOHKwVgD
aHB28d7fo2+8n/YjnR6T9yGSowxVK5jXpdswntwAWUCsM5g+6eKSnoxW0VD6fmgz
Y7qeaeKYuaO72IaZRzVW/qL+kDO/v85zDLmHxfKFmr9xf/FpiSBMR2TWMFVa8jms
RK5iDI2/hbIsUwElG6TsT/n8W3ZBktS/7TfAb3BFZDmeb4Aa2POw8lyx6j6Yo9F8
I6QI3uLfSVKV6CLeKMIql1708yOThYqwehAG9C1UwWW1rHkbYM4Kbfq9IDUNXAif
qHWqJpitriJPCMMd2vQRxTJZtJOUh/W9dou49R1Tc9LpGJ3gxetW+4pLczRbYhhP
mr4h9uo+xwznOEkR2+I7wGEB0G559nnufM4EcYijv8ZlSy9R92d1BkSAmH4fdyOz
ufASEVRf7raHHH4L1QC813q22+ARzNvRVaVahigEG6fySNOWkEmMNXmfN4KQk6LJ
QD/jAqeT2UMcfDVPiWp1Kf1jkrVr+Tan4XvSxv+a3tIjZso4mVDdIOZSzNciR+ri
UGtcywDYP+KWjC9phQi1DByK/dmIPdic/hLkSCCWdLPX+hHav9gmiIDeRRatHJMi
YXdeSOlG6wcJ9Pp/6zo+9Rk5Uc5+Fo3f1AeYszoPAIAd6NfUV3nQ0+HFVz8xYghc
pp8/9jIHkJPL2+dJBl+pxR1aIecPKuTFZMyxoXrLjxZuAmr5ZpIJNdTTH6FBpYuN
oswzXInkpi2vFF60wTujVmQUJ75rBW9nosA0dmPKjRKoV0iVJYVjqP/R7XDAiFtm
yk9efokBwztxKbokNVNTiQZ/0dRXtPSsBX1FauHAjvuye4V41BYEiw3E0ru4HqWq
vBGLt/gMhMOwoUVezzWy6xScta4MJ36mPUuvNCz7OeQWsP8fVv/+fC57ar4VvAKf
2tcBhhV1SRyD+2fXBCILokqA83Q48w9KY3En8uHWLaD68D13AhaTQ0ptkWfeV3Cz
DBSufTgdnJFQx3DmpIuP5oxydkDWjsk98tmj5MDdSZMVeoZT9SnAbPD3kyxCtRC5
75WLsmqyivOuWENBAQdoNsfgggv/OEtf/enI5+sBMy/ujlKNMzspapfEVe/j1IJc
nCFzt91AD037OEg2mtGrNCFxYTpq+H/Q0qXMlRvC92JAp3OWDSSsH0J3M37MprBJ
3PKRY7J1iVT7DtY8CrVsvDTNQwgUwxOl/yKIipZwE7BJFYBn4c1RERf1NNIAuYPz
OwpHsAhTWKW+nmhYTd+7dQhsPC5+dWfkF+jt/h7PKFy05Cqu/fTmQVVl3KhXLGSI
rZUMriPY4li3x92HlVWfaFZ67aAgve35JNeX5cMMKUNdbxzcwLbRa9udVzN/zrFG
T5s+Vypj8LP52D+D7hdkilYepcuppLufBzdWiMI/RvRP3UYc1IbtJdQ/h+QvzTSM
hJ20MmwSyz+uKf7Hzg57iDDyyl+0xUVlvW6H0MMpnrWqHxCOqnpCiKHt2PuVvsdd
n/aRrAb6OfCDPDPMVZCn8+R0BCcfzcyh+QFDcAMGAYMkV5aTtLs1MZkUbNL4IBuM
pXYapELYhwSSM47YPZLtjkZawM0FjSdMzn3jHJXa3TA2fakBCFMqKbO2DyFRkmvA
B/f1fBVJAIbvy0iViH0Xg05Bm3SzfUaPI7YN9fJMJBZ6d4IwYwLAx1hYPVGNzF99
6FSQ9AJTilAvGl4/EPqnC1KOwyDFxzQIFNeCbn4biKKEz8o51nwuxfcfPcE8yKpK
ta+9IHxQvntnN//1kwOK1zK6D+oIFHGEx8chRM9kxc9NJY2R5t/zwi1WTLKJr23Z
/BXEPJc02xlW66j23s7rs55adzppj0qBzR2A1YulXAxoQ62dACsr+C486BPKzttE
FAwLIHu5yEHI8P94HRbqu+W1c4zD4R1n7WHGL0dUyjGuZ4zAoBRZAsON2CE+Fctj
k2s98Z9kte3drEDoXh53fMHUVuFSONProVCtp62ZzVjmzftjQl+9kbSd0o8G5bXj
fETh31l7Ye9FR3DG5mEjayx9wjiSd04a+Te3xFjk2Ek9dxqnAo4i7PqV0ZpM4R3z
LsyLPfR3AlPkyFNYSx/bA91QRl2InqO4gSBOdUCY117vLIF6Owo26oDXkR79e16I
r3Jr3M+rdTtsH7ZxjmYUnihBIHfAwRQUOGZNjGyf3wfIxxPSHekLmXwavdYBIpVY
aOe6W+pJNHylm9wb9mZHnEFe8/I1x60iuil25OPy3whWqbZyHEPi6ZF4T1+MBzii
0O+uFpnpsJnx56CyfaOSmhx+VDCQHw5TqFNbCJHTFwwETDEzXb3VDVYdjo95gP0w
hAwaZypefZX8fzWjkytGK5Gkt0HBvZWGrrSk0bKIpYOz0IMyrUTE7V+9ivy62emd
nagnU6Ad8GDz8euVGpe+qIN4IrmNXi9MTKIhK7jHzc1qQpOaL9xFNjgoBdXdZvQw
WxjiApxREYegTlfmAfqbevHtzO7W5rQtaeUwfL8Ym3PB0JQBFOsIsuq7RU07ERY+
dR02lgJ0eJfxfopE5DyDPLglYtxWlVCe9+Hq/Ua2hZQqhtFfNasbWRJI7rZwhRoV
YgjAdrJYO9nMi0puFFUJRZ8EoMhmw/o9IZJNKF00kUL0fEfWCF6fhkXgyJfmJYn8
MGVfA+jmXpqE/hyNVmew2GW9xmuO4KXJkT/CgXNLVjHaidcYsLTDPdxwyVVv4IA/
3mM004I5yFS6xwD4CLHm72HfQ4B2/VTlNstaJJpfsjCmuSpsOFVtmVIlyjEcXvUn
T7mttIV2YKAYF7ZsZ3mqOcWALjKXOQBVARoGY1/BlDvuw6LVbKGZNd3zElJcSL3A
YWclCDI5dp/1oJq+NGOVO+yqMX8nLGFkojsrPyYrnIih+NMhia/YZhOtJj7+EqeR
fMv6S7zTBnlJuFBHURdzV0N4cxGqVZy0rwuMDvW+VsgS0Ejj6955/ClC5nTM6w8+
kgp46acNxwNDel+S/sJPn6pHGwOeuhiFIiTR/5clMox68yE3KCZWiYOjaoUtyBbk
eFKjlkHwZrowzoI5mCDP0AhrZbYxVdG0qGu4QBDCyxyhItmr95gU1bankfkaWcIT
0S4+1evbp5gNR6V2qoE3QWhp1FKK82kEMooWiy/rQ7vMmvQEWRc6huNGEXU6u9/U
37h1zZ56Ri6UD8OI5RlC7i4Opf4p8tG+xKelbeU+U1hxq8fRzHXqjKjsdja2Xcnr
sruW0E8mt8s+yptYPNH5zxzys0HNv7x23FmDq9gxJ6BKQG+1t6xZU9bEuQoXi/fS
yWmc9fUJfcaCkZlEsnOv3d/8D+JQCcOmFFYA7ZiHGpVlBsUOmrNEO/hVgybc6pEI
mWU4GLzlh2VmZn5BAjHaLYuz8gRuaWSkQRJWdOIJcISP9RRzc1b9N33OXB5YhgTe
VRNQEh8pdm2yFXuUfYFt8MKg36FbaGdkmvQwlguwOY/ac5MDqfSJYIAykht5MyW8
1BpH6N0mtKSBVhwuiB+gZKywY1p1n8GwQAfjS/W1ViQ+Gdb0owlEEaSXNpzNxnG3
fev17MmI50lMpRwYYX4GQs/OjtlZ90QfDzhCoswGyujDcgZuQMrdAVsXgNN4chzL
fJLfNWoiLVXfrj3D4mT22FHL2tb8IvPluMqibHy3QHznKL+vRYSMX3Ii0+G+IDDm
A4miOfS6JL7f4MWABnSO/yg65iyJozjSudXcasjnf835nrsNyI3+Ak6tPLEigeNV
/GIqzMenrSTwTyOK46vAN63LgUKouH++t6npcOwSa26TA+CaEDuk2LcDot5XMXZd
/cMMb4Ko+9SrNYGrT+sut+7Eyqu8f15Kj/lzNqZGY+7F3HZobRkpFI0yPFaBTu06
h0ZTTRatbjSbzBCiZFkwaz4bkyBT5pfrsNMpSIoP7z7F8ZRP26l/TVWdkOgAgkiF
OO5cjJ4J60/wmyISJIJ5c0mwl6CqP/5cqUEHOqdXzrRqdE4tgGg8G8uMJTUqweWH
PPoAKQQzGMsJHM96L6OveRqF6myekyFGz9PLPIbO5et263boEJHRVId0CiZCuJZc
1hezAf6t/MEm6AdwV7ybBFr8savgZYe6sAWKfiUHGc7YeqxMjg0X1q4NTd09+87Q
Kiojg4C2YmDhHxTPxXU7XURiLOjzY1+t32hTP3tzSvmpqTJUmHo1QVj7N2teqGT5
9lxIBbl3hMiNl48YzFdHT2ZgeQau08EZoabrgY7falMndw+LxDQj2smvNwO+XpoA
W226vOeWt3fqIxGy2f4y+vCJ2m9xXDBON2oelRBP7N3vmHK7rIgo7I7jQUEB+kSC
jW7z2r0abRdK1zxBtSxCzN3tFMTylCwrNygnRM8F1ADAKKZ7h7X2byqpVCkQGECQ
BsxkuX8ja+STasVUJhEoApHaTSz2i9vIc/NAHpe6Rco9fQab6SLtVhP+CDLs2W2/
EfAwHWVp81ggHiw0wUoBTtL+XccF0d5waAWI/GxuJQGL88bZ4o2Ay/1mWYXuBGmo
CB2Wfyco9/8We1tTQOCVbQaJqtUFzUGoeHLkVF5JwnJbJX/JWAcPaKMmMJ9+liTc
9sK+rR1GvJP4q7BMFV/BQJ1aXKOyadiD+ZK3W2FU5oAY992AMpl0R/HV/uJYRJgB
GeHik1JcZBEs4Ic0pFCV2peROhHxFcEiodAVcWX8lIWdiG1ndPu9+b/jZtRy9Edd
LB3M9xPZftEQtu4fRmzK+o3qd0lte4ArSenNjx4fiSClY2jxGVUll/D/hvODwxwQ
P3VfbTgdAnbgsRgalKlnJL5Iz24UvqfVuFBnY/85F1zVa7NZLpVZiMwxOdQ8aeBL
+0WF6zzYUD0fEjvI95ypMCmP8MByxI53yC0aWlLOhtW9OJY6rQkn2LXvN4Vs5Hlw
rrHLI97yehT9Z8N+k51jgMPlpYapE2Fffg6iKEkkiXhXAEDLek6iZmLEOO1pePdd
Nog8UcQwLsx/nsIWavtrpDzXVg/QbX6fuJFWZNw71SHyqvdn4xQRSDMrBR6Y9EI2
WxJQnIEYVJIVij99vKUTOke13loPpZodFhBXECe5TvjjzviJ91qq1fylpHz1EQlY
kAAfo+qk/4OUIT3FqBZgfu/3OoRDufS4UtFVX/VkKJ+TiyiHCbcmTIwLsscbtg9F
Jy8EuJps3kqnUAhZR6aX+tYVB2gWLHQXDy+oMNdNMLGMNheJLiHtRAZGqMu04ooO
hbhKf4eCgeEE1Rq1mHAuVgR9DPDAXl8N+7WvWnlDqUnhRIhqZWAH1exFlPii9Bb4
rV+7lW3ovccBemdAwOfo8m32UDzuC6AV/9FHUChcY1ATcJ3GLyo7wK6Fw1PLZCVF
WAXsxHkSajwG7qk5LcbR/HH1ltKLxOCUROwGkpFAL98P4aOR9RFzwl+cVbGvA/3a
zehiRVDGvFoi55fLYY2DvNyFYmRCQJaFT5PSeDWYm/ErR3jD+DitRPwyCOpU+4hi
bUiE5oeUWK8WT+wY3mlNtx06EioK13BF1rawSPkrGTDFASVJKbHbCRd0pQaoYUNn
XxOMWPa9CPr20a/R4QN/DTEysCpQel9WeDMpcJtrGtdDGMrmzOmvCG/POdzvtvy+
e8j+FXUzLSWQEw8uHAzOi9tE3Rdv7qFM4fL1RUHVeAgDOU/Rj5NATcPgkuZdG5GZ
SFIX3UTgRIVltJnv8Vk3Bwsahs/B7HZpv1K+fEAfR4Linq29sC0HjjffGv07tFgi
DqDuVx6sCvTEgKbDArdLhb5v4ROiOM266KtcRNvPE8GyxkxokaAZPXJzLGMunQyK
21SEUbpM2q92Jc6jwog4JDkb4gKJCC8YNRYj8L10je1j6l5ZdPZEo45E1IFD1DHf
SjfVuC1GdWLh6Mp8brA9E3aZ1t4YrhtCCaewkDnv7NoOBFgD7BXy83WR4qCrzTgg
Bs71V/Dcr6peICTVutyVIWD9Ps0WFa1GXjWuQr5e6lRmGsBPWABh+zc1C1Yvtydg
5gZFBC91ukQsOWB4VEn7h0txfH9sBsg48dwTFjK2LiHE1qsrJXI0wy901kq3yJkE
DOJU5YeO7Ja4F+TUwy+Q2ufB6eZttAt/J6NrvL7N53lhO2pytlbVifEQbchIKbX9
SgL5EhO1mewAoju0H59G6YjQaHtAjZ+HvEF1nNH/H7GahDuh1Acm4qqQ6VmFvpQT
p39WNMJGUgu3k+n7jY6B7df8CJopK1+Jy9TV3mnUirUSEBgrq8cGQzPLGVsIlbLg
u8C3Hy7mZM6pLtpbPjxuDY03mF/dOZy7d/QQEZOxibRv0JDcbWRqHX6FCRs0FJTy
5q2AeFAD2Pxse0O9UGxqr+wV+C9GAZNnkP3fqq2B4dxd1oyPAvtK0aHivpWsxAF8
VjwMnQdv0h58s1HR2M65OaDWZOCMEqC9C+XIU7UBmJ4cVL/NknyjIcxZLH4V5Edm
ojEvlhuapxl0bDYb3OkiEPcYHSkrGt88hSYWcN6oTXaQMHAFQxK+WTs6+NKXM2Dq
PD97k3Cr1rmpScEnf2PFog+k+jhP+z1hdLF3u5FMKaA538HmMIgvFqIoT/l/bk/o
cR6g3E0NC9jgo7OIgZbXNKAQpXsQCc6e352RUIqTbWPCez5jGHWWA2nwwKfUjXe7
CX0eHLJpqZg05TJ1SlhxzXHM3IjLSDw6wW7hvatYFsmQIKWcwmqCklXddOWynsI/
uolJfhAadB+jKY1PWCtLiV1NWLEOddlOFIGuONRagwN/1+aCmhehkslDRwKEpkPC
qlJDSAo1OOUpYy9Esm9nVnF0g2TbzjlIOcMoS9mgC7kGdLV8cC6/WTizT68YVG5J
g6pyBdJVYsMxqQw4TP3FaXiTGg7ik5MiGlpEruxmyPch0F4diltbFfXyn95wGWKr
9SFU3qZJq6938157VC9vwr5A3CV/KwaF+F05fUJXmBgdSvzJOCpPsTt0HuklGolZ
fX9pUxPkjJK7nxjXXUxBqxOvtmd/2OgJYTeTpURkEMa83+Pcjn3IN4NidprD1eNq
RTuGRR/uwHRtgEVBJpKfdHBDF82dghpGKtmQ8uTAN6iSHa4HMeYW+YAWaDIM3Eey
ZGhmKS+sA+stf9u5Fc5boRlUvg+IJYBFezaY0D2DsY/1plQ2CRvC6mw0ioxS7Uvn
tzXfSLbbFwqtYL22j1JMfC45kqMvyPrgpWiqb+hc11iVj9emAMdDQFjiqNbOumnG
vnKSW3rCnrsc7cj9YGmGm03KYDjEPd8ZZww0itx5Jm1q0uk8Pv9o71uN+OC98UgK
VyC0L80h8NUDHytztPpCVQYSVbowv8ZVB2ExtnXUnXoexvHUdtQMdob8hjNthDZc
cjHufvbzAM7FI7lthdYjik+IytNJb6H2q1dOYpZKd9/y7n5MkgTbNFkOG3X09y/2
gp5WacJxA4u0LcgqJDcqp4ipfTV9aHobEzcVrMXJ3WeU9nMmC+PXoH1qvD3MnQd9
189L++AfkjQZM8O5UCumyqvlOPs9pn4OskTjT7U4/q9/lYe+yqchuAinNOsL4FIK
0qqQy+r/+FtIOaoZFsfPuKVew4yIj/U9tUzXI0aeWGUIsAQ06FR4Kwk0+iuO6kgX
hWXfOO+8jerY+cQ7FYq4XF8FpV3nM84pEu4TX1MBFMYMwJAxV/8eoQn+bH1imJPR
lteBXSBUm4SUXdrImiZL/19xuwdOpkQJ4n0oBz6C0a5rd3o/1d2bjjzSKt8ncY6C
Rtfh6pIn/la9yYEC9ZW2Cc/nZQWovyLTA4wfv2yTZ/CFH35aER+TjRIBIfIHmIZl
S8MKyEBXflLESsnlW/cumKZaCy2qnsQmysRxUBO++ghVVmEyeWMWtevyjU28V6Zz
yK21pwIVMSIVQ0idlu6XhaBmeTsKa1dXDOQ17HTovDmUg40TjVpF6Ub5d54cGHb8
yfnT7v5goy+npb3TSc0CFiu1SYD1bDVCDIVvzmkEfNeJb8ioMn/NDkHLytlXGE6g
ToWeC6q42s77zif3Z+8ptvCsiUVALjwf8/GvzktzbupaIZQPjJkgQba7pjK1dp0X
FTFQ8pDRqgD5ZRM3ZNp/NHQFn1pJhE5Kle5vzhDCISE1mFCwYkcnZmiFiR/hmRc8
OC1hmbNbMdVmVkk6uSRfIkdP61Py5EihPVj2H86bfE2VUiCzbSsqqixSHNhUW9kg
4fgkAHeowbtBGLp+bm0WvFW3y8dCde/o6rigCL8HaSAZr7rUNzOqAxI1xWPwcHTM
GSjD3RQJyGGEaHWatdtfWvAnPhj2byz/08T4EpDJzWiETBOc9ybY0hHX0rInoafs
h9gayhhQVpPxjlAWSmIcxpPpcLeG/wawnOgXjgBr8bcNq0nbcxYlRljcdtoMu26z
XBl8vbiFNZKHwUhhY0hqXROiIkDSq8K3zAXZRuppzPwCUhhVxko4hdTru+YWoNWs
WkxPvGvSpMR4HwyZi2il04SxLx83qWErfHEVXgXOhAlXoll6LUUZSlfbUA8H06gW
2z/ArxM74N2NDUoF6IlrhO4cxNB80WDi0wd3UZMCC1MmLdlsKSECiiXdgVPzoC0A
mmNyymSc5E3wdILRmiqZz/+mGga6pPZcGCfE50aSdK4rCF0qJjPavRtjBFxER6wI
ho19Fa6v1ix1HDAoXGLcy8quuwSNc8VnnC6PL+hQ4F2aBPEC1zWf2LRCv+oOcV7l
QshJcuOMxCipDPN7n+vI59vaApJLU1jmI98JSMsAXApdy9qDlxcWqfydDXFw81aP
GQ9gJY5dZHrulceVvYF0MvgAlVNHwoxdd8xK1uehwzwcwFinzkwZuT0SzveAlg8R
Q92EONfA6gZ/s+bhgl0zR15R//w4eQ8wuFwN96WESQB9AJGAtzQMn/L+J0Sf06kr
Rmzv6nEZyDE+dAryPyUDlF1ijbeUkXltcIkxKQftm1/1+UrGSu3p+UtySaBemU/0
W0EG75Mw+1iHg8E4oXQ0czdO6K6txf/8khnZimKjr9X3pfVxG0qsG+k8uAYw8oob
W06MCi3ABhEX5rGdHC7ZTRWhjFNrEz1BPzxgQIdUanVdO8zyGbYjhOceon1yT1yL
UWWbHH6raCPvKMgwWytcSrLGD/8C2fRAkSa2M1csoNndkyhTdJh71rQq48xzeXTo
larCdjgGmokWsf0n330NNmtJ6jlu9WAfm67QrHjIkXbNLn23mzWqI/kTi+ayvNrv
9HNZN7kvXjy3zFC2GDlXsoeD3rvf7vcui5bh+SqBCffHAaQ3+GAQonDV6C6QUikn
BgSIWmf5HHv6LV6F4ep1KSy0GQN8HX89Xegd63AZRXLC+PR67XZLgg0FJOI9nDN6
YXIMDTDeQ21IJHqRmygluGVkjjucPIpNy9Hg2cigpyeB7ZC3ZoxLwMcgY8U3SVl9
AkmhLAlHH18HX/nhehko8z4J4FVJybL7RPsHzKYaIF1Ug4vlKmRMhKxlKyOOWavU
6VCEGpREvuz5YTh3cIVLun94pQ+YGPxBdaePKBpkuFO72O0/GlCDm+/drARWgFu3
pNCO/Rr34yzPI/VTGTmtCuC6S9aq/uNtMS/4x2LLOCkWQjFsMeohWfTODIedLFxp
DX9ZtLBmafo+IxyDvcQm6uwsMeUmuAE6OZ2cUxSAMl5EL2j+ZGTFFbyA60a//thJ
He+YH9clOfgH5S1bNy+f04v5Y/xsxrOkkF9eX5dXsCm2eGajdxJPtT6rogroHvkx
A7InZo/X0U8i0DqNSRCoq1/7Mc5HiagYDrTdeN/nbKJDLpsdFayUcXZGJuNu9Czx
ITd4+Ao7HCk1U/LsCFdmlsGdm0scQjv6Ax6EXgtaJ8oJASmRV4BtJjcFds3q1KlR
sYfvovVMybdvS+g1DYH03nGV2gZv+Nnsd0TrUxj+9ZmtCY+8QsMeT7cHcC+pP/wk
//hD/9WNd2WaS6+7kqU3vXp6CkNak+u30GgB3q/jhuaGpUYRtAq/1AgBpkAg6jHo
vqzytYoHJacjriLwcoUEn0hB44qCp25tCREyrMo0+jae7TfRQY6k3bCE4EhZepdv
yjJ+Pyp3uJ1g5a6cVnohG+Uq1nMex4B5a4T/Hdxj8g0Ua2O/K889aCa30ZVq0y3z
sVb5ErVrlQHatY6BAD108Cy7VE7kxlWEaE8nD4aVA5VJWzvOkpKcamUNnWKkWSVf
UNjeoS34jiXU6opYrY/KhzjBXOdL1U7UXoeFGqls4LzpENYKzS1Hj0XklfNpVdqj
KEF8J8VhufmwJU00cQ2bcC4Fk0H7oJcPbht6JQr5FUG+4xB/lOKPIw4gUjhc/03M
wyIApc2IQ86GftNXcGZAM3EqIEZCZ7y9DTpi30xvVvyi3O5OwUjbho24tzCM89oN
RS+qdQBOpdxU13cblNw/pDfdk+dFNsYWo6k7CW58h7wstph/h49FPoULl6AaAT37
L+Kynlemef0XwZm4zr/PhBPVs2EAMy7MMKyPF3xOCxr6wKwbu3JfgbbGEDKXkdvI
6hmj576gDy6bGHGnOE67Giij7KmSXaI9NanppFDg7c9gF6Pd6QcevbHZmlpUQSYk
sZ1lQGcSqMSTzMJZP0m5YiiEAQ6Pjj6SOTSQ2S4cTR4DlcflTHaigCzaeA+7nucL
URrtpqfAsb+WIbg7cEZz5EBA7yx5r7h8nnmZgZw7Q/sAoP9I4NDGQHhw66tZ+ZhQ
SysOxNh9G6cHMckoyLcb8wI25YN0Wqx60xaeMCJmh4GQu0GnbkKWRASft6gCorUP
/AzpYhf27F8jbiEi4qdFqP/5L67HhRW1/rcPj/54VcBbckXRh5o8PORL7J4OwiY8
ubWuGHslH+dy1tJwPyeFvwpBBaox+7wn0Fd68ExKPR7ZhdG+CJG7bGYpWQbnh1Kg
YeO35K28aOMB09neYv6xjT+2DKIf/twjvRqQbQur4DUptqPyfThcx4K64WCqGGAN
W+qK8mY4vrZAelTFVFMmcy7PUFcDk3hhLP5Mq+7sUPb1yR96JI7SNsvTewlVL40H
mcJ26TwAXlNHI1OvjWct2oNynZ65stio7Uij0qgmOE6aRnwQFGAxB41y6g9Z+pzD
FfaCLR2nXMyQFRar9JaehoVAysteLY27fygoXppEze3IeXHRVP3ZlDwo//k0aSYX
xNPcEcSfE7ZOL7Cd8Ogn/I3HsUbNMrKJjgLQt+ujR1NuaO+kia06Mp5GPhEPOywb
TFdgjdHaixJeCi+kLAcNj6WwzcUxKuIKbN8ANH7QUtFrQgfpuzpG/dpimbpRISJb
C1j2v3PtVKWrnCFUoRHwusTgeReK8m+K7FbFWilu82H8QTbl1EItXbdvcNrkfX+T
8JUWT2FD/AZFcyUrYfYR4Ri/gT/e0qcXh4m6WTboAyRj3jpbYPBupNX3QehSeZqa
nYpG7TEXEZOTHnLqdbNBpeuwPGYjotn5tKPuFLSUTJmcQ5xaODe58b0C6peEU3mK
ruCFvnsDiZefTkvVMyExhhUFFcP5IKlUpExP3FqO+50hV0V+niddKwvi7OnMJuOU
qemwla+hIi6/eycPystqSaMdDwPqSYdBE1/l+ES59yX3La3GbMz02QBQD5iM92SD
VXuJVeRwDnZV4K8GBogIRfg21F9dy19H++MqZQRNLvJCBcz4N4O+IUDQxQcrdxXP
tNWEnCSAptvQ2rTnuExA23r8Tj4RPFidbrjxGRQ7aeqo/mLrLBiKIDOjhXGQl+ks
BHSyS3CLaCxuIAZDT/UqHMhr1oyMFKZc5alhQKWlaT3pY2zLhW/Vy+5ZF/4bXWPe
SfdlhQm/tiIHeT9yxsxkXdn0KSD3mVvI6V3jOS0G7tSDnX2NKHwcp01IBrIVKLlx
M6umV3Jq4BDNB8FmkvQ0zXWanU60/uGbeQuE6emf/d9yEwTe4NDsyDV0vq5LYZP1
pCA2ktUv+vVuRQptTXgRiyX6JQo7lCZQcYL7ivLmrKQkW4pHkED8H4fwc7J8J13s
x0VQihABuWmM+qdSmMjoWse3Ah3PUZJgtn4M7x8/UYeVaKZRUKWO9WcUjp0JKdrf
nRZwL/E3mXAdaxaqKH+An2eb1s8u7IOinPvUzTCfjrxTfXRanm7iRuxVchv7/4bK
3kFrGyOQ2hUfj5ftVnvavqLpnXjz09zYVjNxDrSAUQUi8oxOCbiElcI31Ho/jido
MRMp8dHxGzKHLdxuQo0qE9PQJZNZ4js0TTUj7hhfwYV3uL3CA5O/9RVy2VYOKxVv
u4rVv6P/7AK45sja7lbV+5fw0QqQlKBmRjeiavZOJgobo70t2J8xR0KKShZYp21O
CewUSvB1qNSnWConyY4SWlF3Ijw76o8o5EFDCp/uz6PnTrLThanll+UnkwJPQ9FF
uG6ljP7LKp8BnWlMbRE+ntIGVBFrO1qjdOqLrcOF93eaBhewoRK4dMe6j3Hjub5A
wTwo156yUyX4RVVsiHUyPOlVDjDDqYFv0PCRIvVI4C4RVX3GJ+dU7rHUYsPGOuzU
09xnvZ1Bt0yEEfrNaY/iuhYNLcPxDZBuxi/RnT43pjMOMHczsZhGXxjSgzp9s/Nl
QbURIuDR1oj0rBh4BOEoXWXo8lURKhNcYMMaq5SjMHEWD10i2ZiZB9mbmXhCBXd2
rF+Xx+HSO7Yq/iU2fgUJrn55rcymgRqHmRB75IEabUAMCdpaR4Skm1zE+Kt2tchJ
Ck93sXIaRuH5eAsLuMbbpqAicKC5w3q0SRf3OD/IBt3ojTAVo6wzqBrdgvOMWkGy
0pzYSakKjiJyTPWe6lQ6fz6SIcmJeBDpnkMH1/hUMoPImdRVkd0Q/bCaCUvjkOcQ
ER60lPnFvlGg7iP6UvwDIULQHIARSZUg8M2vsJHFRhfB+s/tPSO6kkV8z9WRicCT
w4JEMvc+b/4jTqrkJUAEZMKX26XJyQIscFfSnBpsWFEYQ6CH1ci4R7zryEVEqnpn
VSsN6hzRtrDtUzuaeDaS0ad3VzWe7uT2WsJ9y2XqkqMs9GIzPuGlC6aZYeGRrnBK
qcQwWixo1NHb11IHuJWOcOIsaStKLhVwp7ZrtErcHo0JRc82R7N1vzHfz0/cLorK
e6LGT9t0TrJ4joHA4tM+I0EUgGVrkDPklUWPqXpqBiqFuTUL5Axv1vWDahSLD3uA
NDNJKwgu/nDCn8NcU7cY5kUi7eLeTiKpj1fCBm0tPbaYqs4g4KnOSxAu4Bu4pn9N
1Jp4zxGHsfCdWFIp4vlvbitT+Qb4v5MtqcjZGtH1/MLe48b8KTaoEFA7IaGpqu1K
Zjb4+2Ue4Mb6Psvoj2o5jDfnDOADzJggMH8EcF0jf353hJJ+YuM1FL7SmKqgypuy
+Maw5U4VQ7SEEyixgPn1S2Do02NXZOIN2LV2AoVdoYbJPaQoEBo5U4iRBQsqiEBh
/FkoZQXSOd6lnMZhAXGx0S+6iP6Hd7RweHV9EiDFresJTvTgwVzaXkzHTJrhnhGB
S7U9o2025nxd3lMRpqkMwWp8eIAvNZVwPBj1pXUuwL8cwsAcdTHkAqNh/Djg7dcB
1BSXexheQGOrU1sZ2r42W/2+7nvSDngjjyQ/pyB0KpWtsu/q7XeYGIbLt+m/slR2
ByzU4uXmSN9d1eF7KU/gbL07h3IBD7RkoQ2R73DpmfCO0ywGJIV+qYNRr6Bgsf4P
Y/dgZS7iLEG7WFa0ArfCHWrkHVciijugiMpIOFPDtQtN7F7DcO/q1F4ugdMUQiOK
/auLGEs0tE5tWHWAMAZaQTDgZ7xbDYyPVZCyZtude7W1D6I+7+a05QH6YhzYWFQw
GxOqU9XhsrwClZjINOvaRxADSSi0rI1SyLdhqlXIKLnbDRMZcVhRIwJ37f+ZShVK
3qgeTKb+j5fKMM6zyrkJv/tETWjN5xgzceKbOIm5nrd4jj3JwBJmsm1/LU/W/6jd
v2cTQAyvPwzBmEcGND8JgMe03YdjafIMxHT9p+Mly9SASfPwgguFu2c1+UQ5H0Ho
6eepdIW8a4NHJi4bFMCMTO+6endqjd7z/KVEj7cEsUqe0Qp42tjHFTZyA/zkGHBL
80HQt1ZqP8f6dGCQwGIn2Q7ixLrDohlf9OCfY36wQqNo1C8oPb0r1TdvxFOMTJms
YFRIRP9pTTmjk5LU6MQj6ZhUT/0e7+3o9loBWwGdRHdK6nA96aJVgvZbxSZaWQUD
UbonLXnwRqW4MrnoOetSpSddI13Aiyvgw8UVGT0dSsug14J7i3DvZurTJgVmkLdy
7wIuRCP3Qy11aI5YBr3YBP27UfwQ6AEy2dWkNazmXVrT6cxN71euoyRAHTPv/WhP
WXdG03fiXJU9mVqDEd7EDTjZaObE/5IHmHu3hr4pgBlQUMeif1X31cHRZSuRMWpe
zVFMCNQBrqr1VXIktePbem6eTxg5OjHKudqAg36c3JDQo92oGH3xYLzfwRBTkphu
f8y4/aacfEJZM3V1ZI5oD27Ek4ispoCQU+gxbtg858FCnAXtQ9rComJmuufgAGzM
4idSmrdPlPZ8V1DRWxlIP6Iu9C+O/NgewgJzM4MpTq3Q3n1XhlLSB2Uoem0vuUcy
X9zKK4T4GRsKZYhipnOg55iNiDbXpP7LGAZIUK8aduTEGEX9vmQ6QZvuXIlngSes
cJnkmcC1XMol5D4DsImzlWz/SZSKWsk86DtqY4Ivu7/0PJxcjhs+s4TQBJLtVoS1
PZ8/gwfbp4zdBRGidboeQgr03pwt+mYbKx9n5u2/wYF4uNhQaqyTEi5BW8K23f6H
3R5rZZ18YbkBN6r6mCXU0gfy0UKcPclU756bfiERvpp7CNDoDqgHBXQmToYg0zm7
F1h0hC397T5/4T831jaMvL7ACcjH9IhYU+C3eWFmpTw4sqoYdQs7YkAbP3FoIbuR
UXuju8Cfr+hMqFM2nVJKFL5f/EgLxtMSMZr9VGNQq19DzS9m8tgpQXAJyRuuxKwT
E7OqWZNEVk5FCneZ1HYiAXQ7SMSlfuPPWam3izeT13Oro7Y47MaqIjv+GUjRAkSU
UCndRH6clwA1ZypbPGt69O7cDy/gZbFcpw2kP9rqldx70xld2OfF16DLIVZwYy/m
rzvz4fzOWRjRQ03i0U+6thNCnw34/ir9m+Ekll5V9vOoEFb1pTSztQk89AOwEN21
aJwFft1mNjjvnEJoNAwgXXes1TGbpz8V+qmfA6+6Dp9A2/0g0xaUO1oBlNxB770a
QxnWMggvK2WKRaru3bn9mJNIfUWjd4qbXNSMbI3V7sWgjZDBVcmu3Cgn8lUetKfC
TKfzAEcEfzBYvTI3EYD/lsCFVDM/zeTvUNebAjHTSfDS64BgTZQI1G9sK5qpxgQn
mie/j4BP0HF5vGQAiFqX7bseCZb75VtTk2qWkUnkBABAepG4twW9QsPfld0gBSMa
Qt9KHuiW3qXrhtahoYPvUHlHtSjDrKqGSWB15klr4doKqpeSnH40X8Ke3vKs8gWL
MhejxXKTvH8vt2H4pJTAjZlBVnUwhZyLTm/MpsGFrYYdd7W+/Z80RZgghFJ4kqfT
HtT6+64N1Ll5AQ3xCJKlg1PrxM+ymC5S4AXj70egSX2rCUE9CTbjS+DiAR11nOgh
xRopsaReXHy5pwC/tbCgelaZ3uHekk3cC0toL2itx0T3Stgk+7P0DNWyBWKRKRTo
Sj5oja4+PlQIpTh8U0UHmyABa6qz3l0vGp3syMeeaIV+GtP9J7vMJ8pECU+ne+f4
jLv9J9MYk3g/QAhLpnmydPGSH2gRUIB4nV0AkkyDK3I94rUjk+z5czE/yeb/zZdn
6KIILUzZR6AQiKjkNskNGWq9RahTHmUMADT9naA52KbtjYbdKIOnXkAB5wQQg0sC
VriWEUDZj4IiERhcTIoDgL1tX0K6DCd3Um7YslFDl5piuz2qhy6cnY1RGkwn7prF
CVG0U+1evYTsPWDkdy+BnwzENs/qtVvFaxD0Am/1eT/fQRhwD/2pnvfogi8fhwqZ
Yz2duuoiJrNINGKcIe1BAWBHKzHbO2XD3ZifnoAsVhJvZYXZkBBGVRUSSltLcUP8
YQdapenstCIupihxl1jc6R58+SRk8dpSTREgR+KQnF0nf6QOzgAZC0UW/76HhNOq
4Q3lnJh8M6bV55NHbkgA0jDjdbGFYVjHcQfg5ZSez6tPrcx9v7qZLTozR49ezNyl
gb23KBzYE4NYL3DzWUUzm5y6SNWcHbHE8MUPTh9CmVJnJVIwOhTOTj07Xk4amc1G
Oexms4bngNeV2X7ZByWTRjnMLP8Rd11v/e5alF4tY/LLXHrV7+yY/FW0P7wzlv7K
FD+61y+24Wll1PGL4uRTe+BCGuzbOA2iAFdKIvc5rf15iWQYTbR5L4Hc62ntZM3c
pIbPQJBSo2qR2v/J7c840QaV5oDSeBYnZwAZbh/LsdCNTnbtNOE/C55d9gMTDHbK
gyLzNRlPUa6utKZCKtyh15X6gvbnra6lEuCcSrVZmHqtCtkADI6QZuyX9hhZT/uC
m0wtOZetvnnucFgxB4GaA1ePtI6xopu4Xs7PuIFuXFib92bKXFa8zswJfDAKQIXJ
qkZYl87/SbrM6cbThh16dZpTLNKiHTJ6g8cEoKICt8HVkEfTDqintFkaHGvsYJJy
8w6JdBYmAdwz5pre6CBOfiEYk78+JFbEgTbteNte17iWmTt4wenQnpO5Y6bwdV7o
lzIzDlv7/Pk8jUvSfE9tI3BQ5FvOjpqKBenbKJmVK7To5HTDoXTzet7hXTKFWtSB
67y8/vRinluESJ/6D9AoKa12IAD3LTu32qtkSar2p9kS9kzSBp2VkFfAo7KAPLtx
zA40rgf2F988IwWyUO88KsETKXHniiFuRzNOBUZuzM9iJvhCnkaaF022CYfjcIIe
6ZHKnnlyB7DYm1MnDZXCZx3usjiEeknJga/hWShoMi5/9hG7YrxCkmXzvLj4l3N5
N1KrZJ6jKqFkaOMyqDQf/yxFRc6rqVEFzqZMQCjVxCqV6lWK18idVsgXGGJYZQ3q
X7CYfbwooHH82lyhgvLFtLcsJrDs1fIJ0sNCcuHJeCOEV777P/Ty3DlApEJzRXeO
7AoMgP48MVddjGoaeOp0vQ1izpaBLK3k3lINzsUxdFTHcfE3wvBsW8hWoUYyr5Z/
q9DbFUxT5vagOfSRCWsgU3/7AgzD1nqh8lLKGE1wT5d3RIqsXT6mTJJtyummIVxn
1+6G5l09rb6ZSfp0jylOGRbqXfbtZqYPUY8S5F/VX04iZGerVvYLnWzQnKZpGig6
gpMsZ5tzFTFUPTcVFE8KmWobuZ3XRXVX9clcBCMsJsbshuHyJt9qPei3mP/ZNhXt
Tc+1sGwhGUMhz8LZ09zu14IrtV3Pez2fpaTjTjG13X68qRrvAnjTDp7q8V4BkAmR
fyPVjCv4H1H9OX2wM4k4xol4bFGJL5MnrASCr4Y8SQz8ReZ212BfRLYZKgpNuZVl
Vhjpi2s0aafyqJ9cj5cwaST3Ic4+xDnrWv7AMhzeyB0OjSzVR9a8TNYhll3Y97BQ
q4w9tIDMLN6deAjBeGsqocY6ZPtAOElJqdd5CMaaZY7RyuHXjdm7703gI9aQroVS
kPIdpoT5m2U1g0n82l/ZzTNmw99KQ00bcdvvVok8Qbqr4ORHOxElY7wGpTqyfzF7
93R/hbu/jwvlHPXFPPiSu4vmzqK6MZSo9rlPrF9ZKRoRIISz5hi7uiufZrmOnRZY
10CWh6YXkAf4flu5HuG1xrOP/yuVM028ovZQpTOPUAXpXQaAENq9Jskf2Qs/qgSK
LsMfcchWZeGj8EV113hJadV9Sz5W0+OQE/ID5JmRU1JOubNDnJ9Jcwl45yBJcAXH
1Qe13w32S5ezEmMAxcFYBoVt3F7QsyG8zuL+w2wnAQfRNfb9uwXisYqcIHSNI1Et
0ertwBvHB9a9xqQ/tGe3i77Ij1JyJcjhg7HAbn6y0Tzldv46inhZkVStjgIRh/by
ifn6Ti4lKJMsH+Oxt6peJknc4o2XwBSRiM1Eh+vrrUl8bA2NiKOeqvou67sWOWzc
KigIBA3xODTlKOLlrpDC4sWOicLw9Y+vGylN6T49G4/ehmyZx6kp+c8CFKnCNI82
9DqF1J5TF8TQaiopB4psoE4BDgvQ4aAwwNXyH0J+Iu9sxindhvZ6jsZKr5qq6r2N
vJCgc1PHS3sbhVfau7VPX2Ejd29Y9M2c6dWQIsuW5x71jVpHhD09U0nMU6TgpeWK
bBKO4nIG9abEPjypYgQLHGriMye3Yqm1NPNWJBtwVncGPmDXZK5m/tFXz+JNVKad
vHfZNkmenbUpfQ6ZzXeI/3CDXT+GfsrdYJXzQwCjrEHAg0JueQI2H0l0pjaOZi0m
rD65H8VB217cXHpFbBUwBiw+0fzCT1dYE1Td+CN8vdZYAXHJQXK9yYsZJ7LkGH7g
lOSYc/UFzOWudDHtI0jUC9Y2PTJoUQUVBJ9V6npVs/wI0Bp3ucmBrhArClWkGav1
4UeR+xDdP3XA9nwB6Bj09rJrv1ckIBUQZ11TJ9VoK7GKZ9W+vorEfJlpS/Ov4BgX
711Y88ky5EezgvHVzsTh4uMuqk2spRNEceTRNinkkJF6fV/20rgV7V4AIHt91Uji
wirSRRLTVqNpigu1ols1Kq7CVrSqBIrWkE8fhWjk/0/Ovp/veCbelELRVsRkueYn
95lccH4pdIZyzQT/LVHYmA3jkJWS+XUDL6XcD4ALFgqnKaz07y3ITbZ5enidLrAI
s4pgY4T1bsPXsuOE0HKqyQJdRnPW2S4uB5BZxs/z1W4McAxmbD3oKNmmG7dEb8bp
Ayb/xobq0ElvF9PBFzBTrNHr7NndbLrT0x5pNk1T7ryLo3wDdlH7iffWiZlSaDJ+
/AaMfqD2VTep8dr2m/pQiKWZdGSDP9Jxum4Ss+qgsvT5MDlZEJWkJbHMMg4QqTlU
bVoGulwv/ba+bbhsQICHchV8qsz2PhOLB/Vm7uGxrWm8EEF02R6IIoV1UJnci9cM
1NAyjWtUp0wofC/YkhOYMcKbRG68YuHK8iy8OF6kVoOVa7tS4SWvB0pYrK2DY5RY
UgdgO7SwZP4NCJzn58wVmxRume/kKP+OBQn0UhrCtA6UlTkXUtMa0qZ7mbTj4KiQ
V1Kh6JfxoJj9uxPZNAm9KhV0il4SrLtKfffFLmZT7dSMOMujWEiqXMUAsn1h5qCi
8eCWvxsppu236jWB0M6nbeG+52NNRtt05kuri9w8/LP4kcRmaxNRIHI2Bl7+YKpR
NpcVZSTS9OV4Hbk9FJUemiT/YLRje0dJVQZ8eH+szKEfvUlWr0tV8ISwjLrcwZsu
H481tr++prjH6I+OnByesDWNLdXys+hjSMpGsiKGqSCEJITkDvY72SyIMW6WdGQy
FWIoplmYLGjedI5NRjFRtBWZZeeIJmjhy1VJq4kEpzRr0sXaiwPnoZlFL8k855hN
eoZUTlYAOegJ5hNp7+NkNtB+FetR7p4uU76atGYzkrgAeocGRc2OAK4riOOyHEia
m1n50RHNk9nIAwVW16Uwh6QALuE8w6E94rbogn49Ye7d18UUVYU6IBL1tzrLTDje
HRa2R7nuH4ICwFcZZ/vEDsAiMc+3jKpSdgIswx2BCA3AFaE61aQUVvjWIIWjWUCN
3sDJFPT3XCHztNQODISfPRE5sVZhc0csJDIl+7t9BOzCS1izFQdmyMTXs11pxVeB
tt7MS1PSi20ya227toH1bxSMcDcyfHzqKuJz2O22YBllgyEMEUfnFZqq98W2HSQ8
EbAWsuFlCplqEf+Pnbq9kjX2xHDcZZLa8haQ7zeGcLJtdlistuvHCIXwpp+ch14n
ouEvikGvQaEgfAyQM/TiKFpAhzc0Z3XDrZ46nyydlRkhQ6uudmRsCz0ZJhgDAAsc
1RecVyTNGkHH1jPRrSgRS3OI2PfOGdvb8NRH+VMSbJUqnuhAo7MXFggse0uDFIuA
0bc0zoa3dnKmlP6xLMPw5oNgOTQD/V335E6RLnbl34W8W3O7p9rDQqz4WVqFYR89
FONXEzMz7rgZ1SnZRnfKpru/ipxgZ6qa0E37hJK6zXG6oMaTrdRMJeqzW+iFeKjv
LrWUL4YZS9ubqRbBMP9LX5k/HAU1QpZtNaNzfS4p6VApyLT4CZpQXggzQdDtDonT
F9NXCTnRszWY8lnr39RQmTd1K6m+NisZgI3IoJnt1erYhfAooFI4eKYTYIuQ8LsP
GlmJL12xU/DUBLd4LvaLry2PBth939r/F1txF+KohywVUnP8+54i06lGt1uZAqkO
jVWLs/f/44aM0Ec+5QBoKQ2DiDCubIbPFhTrOcXsjH1mMwEUgzyxwsC5nFhD/Cwi
3j7mt1TgcZqiKFDrahc34NZD+IanVFxIn0p8dZzB+qcRpPYLxdIF6b+A/zlJfulf
HNCsk+bYczlu1eX//vGpu9wQXBx+SyM6tmtCDrQNKgnpWP3Qd+1lnoi2XGwSdWIP
N72pmhPNGAgdRlDG1vutjKpY/3jwdl4IGcL6uuDxvxBgi+1IQNsXREsVaUFZEMLE
zNLF9w2mWMxte9hS9JWCIPawqEPYC4hhnb/cmRtNbY5ltyd5Wbr/W3rDCHMSBJuE
DyfHMpkcqJ48eJ9IkGVkXu5lqJbjR6ecLIbucNcFOC/tCtT01AlcyCeVUgsylRRr
1ULJioT2uCyxrYQc1tS/34PlUANnlBKT1SQuXDZL9+B63OMeOL1WN/NgnFf5ya//
hhSrOwmvaJHTqARyxQgg94770JQRCe1PU0ZdsF00i9SXVGods2xLTh8gl5TlET7A
kb5YU4wTNIk8TdrzK2hMS2bh5ocZzN5RG0b4c6Zt0Ib4Oxino15q9tvG/PZnC3VB
gb44wicaLhZfPAshlD65hUPhq2yOUhvZgg62kIY44PLkyLZnZ9hhBNis//mPDQx3
MdLKpaVnrliHKWJMIHDIonAqp6F8CsQ7SqmgFSa5yZxCxpNXwBQg/KTk7iz/FxIp
1SkTfLVxn+0AkjvAoiH/OnHe2m2mi1kc8ViXe+pZZIb/iVnXOX+utNu1N+2xPGeh
vvWp01AxIEGxbvIyhWJCYFmjE2gNYOPHS+Snht8fmsnqUl7QsVqRd1pVbt1HzcdP
ZbC5CpJ+u3KQanPWQmuh9QkxIyfeTupj4rovvLg774Nb0qUYoCgl04BX/6lMwnbG
zwfUsoEuKqiu3whion6G2qWsW99x8ZMjLZLv53Hmdih6I71gJmvwLC32FWuI1WGf
BUmqhZbpBNPcAizPc2voG0xxjgiwTsv1+IHzGXooIZStyObM5XzBbFYa5z20qTqa
m6iuV7zahFy5t1KhRiSK6mWIOM9BCSwzfhnH5kzO820uNrpsgNQz8inHQ/jUbF+7
hZMAvFQtciC3FH3eY/7bdsDtJxaJdD/3f9sqXWN35PzKWuuyfKQtlMNDyMkPU0CB
vVN8hXoANvAQDMKIcUoL5gw7Tg3rmYnI7JcOf1taHjk8vaja2gBua82/JR71mbBd
PwXAXZak8C/ho00krxgyKVJ6R4vKmf0AqALkfWiWQywYrtyLCp6/HcjcQReWwTGk
FpwdlXfi4acS+IM7AlPX5IXyeWWNR/h7ZtiHGuNEDQQgqNelsdHaQqb20Hm+Xa7Z
VUN9yrjZMgEHH+nUs35cVLlIgWwyaemCfGyd0wKb8BJCLPwBBDLNVKwNcTF5Azr+
coO17A+KyLwI95XBCLFTfc16/X/+4/kq1wyuI3fEgvVN3wdk9MNLUwt5mhCdw9qa
MD71Ish78mIg8ZiMZJeuaBrBEQVNtkUF90DP7Wav00wq39Cc4sEUznIu35ibrU8S
sEwJaLxkgXAoRgzcy1Ix8F2HJhNKM4+y0TjY4VlUtt4H5CJSKB4xgcn4GNtzrEXU
YFk6oDnodM8HlyxXOt6EdL769jXQZpXSVQ8+W5y6tuwIBk4C1oTpbIflRNA2bj0L
ZAStq2WqjoLMBMDLrbe05WAmFwVdoLlEXtT+HBFe8alggTmUnw21QBKgpGexOwOY
aj4UIjN6jwkBwIwmW0Dr5JT6bFYnY5fj/5iZ08YM5bFpwNYe7vvtPrDtd3L4/G5Y
fNK8G6ZryuUdr504wFLPEZflB8TTwTx0Oj+V0hKegolsXHnJcOBePSsLfaoU4isL
pANFk4p7BxOTsj1GUmldGpsVB6Wr5/WZV6DCABTUP9NWsvGTnNgpikH718okkacW
Cq88gz4BicewKXAuYqrvcFULvvAM4PQiOcc+PShMj/SX0czuseXAGEh2hcdwT0fI
e5PTppJslphnLIwPDPohmj/oNOHvnaX3/L996fYu/JVRVe9qv32Lg7fOJr9QjENa
RCflfkLto0xW6asS6594jxz0fxORoSAXMgWg4uUptMzrtCmA4lh2K0CmYuMh6wq6
mdskOsFiMh9Lb3DanAzbNgLZNe5uWDwQhlEJ9zdodm68gelnQ/ReDD8bOIG0ZhLD
aa5roqTqbLbwMnQgK4OqusxDJliHRqOVZqvrjK5G0E/VEyJ+7jAiL1BxXJK+0mo+
+KEdXhJPhbOe/w9YKjBYeyyAvS/ep9ixZdH/n32wYrWvzFxy4rgZFXvhjM2r4SkN
CdkuI2LDWgIuCRUf+mINOxrjdR+cvYMLSRIBgTFnCShprqNuEeO8g3amOJsLlk19
sMJc22AYW3d/mkWhjw/DFrTNi93pkzvVg8AncIDQgUCQScwXZLui/VWRyFPQssvf
pHViPKOeeKAxRSpSNG23MGUNupKAyGkZ809EzR6s29qw5ZhHw5wPu3bkxIWFF36y
SSh9ATGLS4PCjnUmWP7Ul40phZnt2FohRJZQ/1XsYRCC1zVcqosAB5a0xcvv5Mq0
ZLsRatUIbXpX6ZYoKdyp6Z0Rnat2dU51DPhwdJpYCOEibmOfk/E3uDPJG36tDfd0
6P5oJ6p4gDNMOh5OJl5zsGHqvl7nqdSCDDMeNek9G4XuL4zQiQrm6vI14C0jlDmM
LDgKLIAN28VRszUiPh+eExOBVc1HbE82XPbnxAj1hhett5wyHs3Fwc3IsMXAWLzW
1qh8k1gwupbFxY309jr48tbQq31KPaCAanuYdqRq9FL8l3y+hWXFWzrnGUeJ1VEa
we6GBCxtVtIdpFx6uJL01nDi9xNEAyDjmfv1SJkeLA8dHUWTtgkfGp/qWwVvnKZK
fX/0jhgLT/pyMBMg0Oy5jpP/kTWzFzKoSC9gyE60F+wotegzScBs59IJRBCXLPND
17Vw3rPe6v+StkErqFFKKhUnGq7zz/Zk8Qhc8ald6g53pYOCAdIVagy7JnnJ2vF7
Zr1hVRuONJhFvwEsqWGpADMZZnjAP8DyvEh+YaboEN8LL8AvFwsW77/uRBL0z3ra
aUFb9/QXkTr88o5euMK1yrc6mncPDoO1Wt+MHcxQyzCL9M21HKo2/i6/4tzc4aH8
hgJ0oVpsn4OhlhbrFOKBWHCFE6sObAANmYkZaxuwE21UOZZC+at8FZrMYEc/u6mF
LBjhuUpiIPmK8oDxSvXny8c/jloX5z+VNztFi0oWAgc3Evqf6jV6alec7sUtmzBj
EO+dcS77qd966oBmLK0mQCeX9OozRrfwc9wmn2URQHXV31hUlkIKUzB4T0RXTPZn
OTiqPbGVQK/AfKScgh1YEB+/2iVHpta5Ot/5/7SdaOpbo4ErnP37D/41caut0/o+
ROfzAMn47gArHx/z29vot+OwSynJxNJhhEBN/dhTxke1BRcuSQx/WHbNzt4jEuPP
1VsLX7ArAC/JkIk3smHqWL9yNMmV93pc5kNHfjxb3z+HfBo4zKvAeWDPN2ZTyZJp
MMPYwCTqxQS/s67R5qkI+o4jVSJ4AZ5U6Gbs39KjgV4unsi7CUxzJqMAv4gGCHa3
8cx5hIWAx/SUaqPePsDNzSpoUpiAUiR/cMBdIAKc3BjM7zob+V2U/q4Uim1U6Use
a3u67oePeCF+INERNdcTKTTYV58NxqBM20eBV2n2eZ17XT9qRAQUfv8uPz7x+jq0
zBiTpuDVsq6895KNrBTl1/vDfuOX9VJJ8jcN6oq/k2N9tz1usiIi/Q5MHFicKC67
wAFG2qL1n2g8JAORAnECtJ+SfYO1V0r43WqKR+Tov4ZKGUWA4XSC+Hj9Zdgn620E
zfXoD37uLQ6KAGvHoJbbRr2Zb5t8XHcqsJruF5dXXIl/NGYuNkbApN8t2QAYLUV2
yQo4dXYfRCdVFSkHz7szHWR3ffLx1armjXcTA4kNcCO67kTgTCOIbLdAjBeDTPYy
KBkpQU633fx2EzFkmjbarAH2lrqSegVQxfDbgBecwi+RxVx0kAlONtCfBCoR/i9o
zm40Y2xh0uxpb24l6MPsP813Na76qmNfI5D+ZQrSZJbtIicnwmu0nw1UO8LF0uh/
CxhcYRgFZYBaIEHELAejRogFgvrFt7D0l+/ILm4ewzwEoSjU6vw58esXFWIGjMK0
gioYp/9tF0d5kWDQF/JjYe/xjBeCtaXB8LyXQJUiFMkRswDRrTN7oVHb82cpTGPZ
N6PhsPbZiV9V2aO+DZJECxvPB5SbMhOLJNNkYlmzAetYW0oMXSyTx7487CUNdM5/
Vo1zMxVURXJCTVtStHaFtSYYzHdNMB6nGtkjJGtJSFqseSqWOe9ujgbk+HwfKqnT
Qj7NpZD6Wuhl22U/yPXGWK1KESKQtmB5/IZi5P+dkGT3lPJKMWyz3z6sIIzciFcw
BNMQgy4B4MewlEKbb9x8QrFzPzG7JaTnE5CDXDzLDe/7bFPCQwDZ9MDHhFVh76Ya
U2Dpq52MNA4B5ctAZwGvhfkdosVXStXWw8NC4K/V5P6/oYC2ZZUKaON6bdUXPHpJ
pgrC2VaDesOMeDQL08j+oqeggVhjHH8qzRaSzqfK+g8ZDfxgQWKkmIlmdvzLQP/I
O3/6zAFOJnH/dvFA7hO2GiEi6ANfkB0K05pxRg/IN+mimBc+Ityp31oqrmcCpYv+
e8l+hsjpazPocJAylsoigUOXjjdEbodVcxoPIuJ+vOmNjxSAMNvwF2sQcfxR3x+P
2H3ys3DSbEuJuyq9avOymR/dAntdVKw3n0ePraguoDNgAa8Jn//jrwMfWsASaoMD
9pHtmi3p9HKEj0Q4MkeVhD9TT2YumCFqoMjzJP1YcrmDq2oAyARnb08DOK1FJSW5
PfdD2R6PVU1BGSpFFiVlsWsYvxU7LodqDaj7m1Jqm2RNNvv1/v80eYxTsGmWLb5A
O6TumrVXavB72oj0KalUifZCZvE71E6QJAm+AVBTu8n5j28q3KARKLPJ6snszlN2
HMVCyUTaXlREgolDjyjMjxNjxK9/cPSfarTuqm9iEbUgAaX9RAlCq1kKo3fuNbS7
2DjqcLkwVsYvxiXJmBbiQcNVs6TTL9CVVGg45byD7mPH0w8TyKSwT56A2DlBwUP1
6Jbj9eUYh1HyvUc18JoAKwZO8bEYOV24ciP30Lj39wQG1m8+0latUjaWGUn1w+Ud
3aehgugVHSmCEkz6GuU9NTHRZqHXXTLtR75yjl8u2v5dZXT+g9tDdGUsTOwtcIJ8
EvLHkoYgm4llCb3LSj8VOBJdxZRPOQFRkKL1MaKyWfwmBnjoJVbSKfJ1YdQYH4pJ
V6X21+Of05jkNNiLJ1FQ+7kCKNzFFNc6KziwR7iDkeK8ow9PfmIbO1020LsP+csv
QNijBBxftdwoQ86p4zdJwJIBoTkOn4sW+4rwEg4jb/XNRHYxr57BXozeQHVuHwmP
tXfQiIpA0PAFJLy4QsdS186dtAOrrVFeRD8ppzz3CA64h85xTqML1dTFvhFEu0Sl
t36y20GCFzHGF/2zhkn658sXpsqbigsR+ERYC+5klFmFY03jzCIwQl6QrQHhE3CC
UfCGHHw1Wn+hOVJPqVBzPjOmMhueu3cOnVzREfYf3hOTCm6Hq2Y+AGFi0Nfoc/gw
D4ziNlNVklXTqFacaeASXU5uyu2AqzLNkzrHGvGBcbQ6X3BjEFHLK65hDZi+/Vni
t7D840eSAVUrq9d/G87X4EHf6y5LTooLngi/QsUWBiXmRdJoYUvamoLay/JiSbej
bJG2YfExXGZFaUgrKW9gX97zWqrCh3RhnquB5DicicEYSl710w6eQQUK2+SBToVY
43H5h/DDif2bODqlyKm7meMrbn7hUb1QbJTj7DfsnSdihe9yXajUacjb1AkvV280
vCYj41zK34ZDz5S02c7CUTFM2lNaJ6Hm9+r7HcVKQmB4BIsTjVR9NuopvZLpDnMo
l0azph7oDazY13qCqa8n/NOZfn7H+K4eURS2P2NpBeFvJPNg+yXxhFnxgAAFAi+/
DFqPKoxVaUL2BM3Me1faIJu46Y2Sm+77qqs4FPkfCPyPJxVl20asVMu74T3IirSx
gQSCjOEj9ByTYbE2HlviMUz2K2zoAoLBfzDuTNRMUprOHrshbgPoHGZdK5u0QRP6
oiE6zjoBqxL/bjVQgpdb7+bYQmUnZnTC/QJtazUTSu/ab41K0PTDaZ+lmYTxo+09
sVyMEBuI4CvHYcVCeJUx/Eje9TPP2ryizbUjVgUFQRZ4xQyS/zMThNR49KwW7Ivi
7Hlv9vGmvznxINUNGuD+J/h47YLRL6OuSrfdwCM+cQxXDYGMf7m2qCEC4+dJeaXD
dAD1z28CQPBfBOZ5tzoe7/ypS/A5J+NVifGnnu3UKR0gxlfJ/5qyoAaKUjI2Fv/j
r0X9Kk545n20D2Lnc+EYMV7W+JSLBUB1NNQA2SFUGrJ4YL/MSQJ0R9zodjbDdl56
X6P6OiiTMihRmNbuyXuhyepceqavJqKCBVo2hoydB8a0JCSjfl/qAPxuxFInmSoc
jvAJB9vKZAXdKmchVMu8/8ZKka9eLRCv1Lr1mEbo4FBAeOPCw56J6jdOVaLfLD98
HxGKBqvhbw2GvhGwvKr/PS77IYl3JNUo9oBEzV4NHgCBVAw5Bi7ZzmwL0vOpLBr0
Rt051ABoertfLTQWnvZPk/0UjcamaJc5De2rL5z8MraOnUtvX9eMd92Wv2yMvBIv
mV0ACjZSWfPyJW0u2B0a9Gsh9EwCInykkJPHT7Xmv03R1mxEJpsSSP1SV6ZbiMke
MbGC2y3LFSHOYrjnPWJ0ox7fOGWlxbEbI62g964Y46HfXYrBFZIHtk2jPR+mdrkx
RwSXP9OvQiAJhCx8q3wQ/+OkxMaV4XioqihE/Ys9EDRGbeVwCwXb+FjRL4txz8lD
F6Ag4gYSeLM7D7lrnLFgUqCn2ewtpIlzdGubj2NCgIAGVrMXc4ArXbXvpYKbjan4
kkJCechPxasxfX8VaYMtc+3bwzEqMhpK4C2HvOb0HO/3qtnPg+Du8Za1l2rQnlty
iCj09nvMZa69pTewBwbyTyYOMC18PYfT0sZdUd9MW7LairlqR/OabFyOvth6aE7n
7jcGgNjKBZxPkSa6OwONfu+ouG8Hi9eYez1Me1K6V6lhoZgPYlWexPwtCfOch+fP
9TMBWwX6DkSY6Uzi+3CiDC5GRZu+cMdLOCoqYj+To4OHr7sWtmckVYk31NTbx6Zk
DamHpLerIqsDD3I1fy5gJco7R2s5GhZmCYB24xsNB6lMzSjy4wjRVnQ6w1SZDlVI
jy1BFToiJKD1JufCWApvmj7fguJ1UxcLX71SJFJPfektQAdU362oj9HMkzaUezfV
Ql5B5GvU3Rt+eaL+HW4+r8SlZO+feVjiZIcnJFuhPtX0FgqNuKHZ1cidhW5PkFsY
WRr2gYnZiJyHXktluUgn/oEfbMQZUUXL4xAEHJy3QNsT00SRyljj0DYHfF/3yUIj
3Ia8OVgxBRqTNVrrGCCART405pxP1kD5rPFldmceyiX/9PAw3I2ro7ZK76y1IAa1
32xA4syX+GstSFH4KyFKaPWX4bkSdx11n4rI0HfHdcsoilkkYlP71r4GuGhdk2xg
YpQTCR1XLIl2QSfTamepNwp1FFGhexlxvySaXT8jT7hfjoReLSTqBJPXB8LZ8NGf
85riYADJcH6OEnec48kf4IVT56QFmsCq3P3HdN/j18fMmjJzZeO2a6hTEXtrJ7oE
pC6kURHSA+sRTBv/jv4d474Mm0omwB9T6gJxweBaw1PBnl/OEoT91pYvU1N/AKSJ
XtSVgI2U2FdbcJU+MFw76wc2zZ/l7lp1Xhy82g+M0wHc63DDcS3pyq659ay+ZUbo
1EhqZ3Lz5XLfrgAmP/aKSQpUMztA82ZiPB9ULkRy9Bi4yRkzN27WMaCVr6aQz36G
gqrjUxX6t5HB7tM4FTtrG3vC/Laul1HOXnJblyVnEeuuwXgtHjzreUoTUUIochDb
jEHJQVpdfT4DF4mkodeqYK8HpULef+QhRcMFu8IHvMO+of5PYADbcr4ZT5pPgpnc
FWUdZ7QoHFVcZUoO3oSFucckMpb/QRsk5HzXNeQwEaV5sJo6z72koE978zDSbvGk
7YlOkV+NIYifJBcKxcqPtf8kEUiSzpDxo48gh8O0dPQ+O3YM7PsW+oFJomQ5auw/
Mk8SlCQvp2Cudgtc4fAdj1NNg98f99NksQHK4PD54TTZsP8HKViDR7m2mVTBnE9h
SlkELgMApnTNp+oVDepGZLwjwq54Y2ag3JHFyEks8xb41kZYs3NAg3tuOcwWjXZ9
bu+HJAi/N7pBIV4nVsVJ8ylgUxpR1pBWDZgtaxvOsvoTiPPMLyRtiaYzy/6tVOCm
Ilr7otc+ZZaJqDOya03tE13og+rEKvxyDbHpltbO33eW4R1RO9QgKu+mco3HY/RI
LHzthzjpoj9L6mNB6owENweBPGS/ILuTfdtx/0j7Z2BGUYxSPeZE5UyYeTI/PPHd
UfmuFP3jO/uRwd61odL1I9q0QRpx8o4tcakXow4rIi6ZxI1kGqk0eqB8y5QSkMND
aLyf1w/TWgZ6s9takXZD+64St6/YoFsLoTosVzc+HsN+4HOh0CPnll1Sr/1S/zY5
dajYwoxJvJNTkkAAxdk4vqbVsWqWetiQA2UIqrJM6OAOrMtQF5hw/Bo0QpLi8vFB
XJJRrFeXcnEWJ4qB8LD4lQK0oc2cZYZndUdM1rJKv2/paiN+U4AeTmNd5Fs6RIwM
tLfFOA2EdHwK4lIXJ8xPkv+2HAriyvHtZgRPAXlsNltZizQzrVLYAWMsDlNjnTKW
LVj2TtKpjLyoV7QNy5936mZSRpz8X+OM1l/3I1GmdQJPrD/jCVy/gCkivhJmWFDI
88wlN/o/EQ6hqZCsPQDyQJnIp5T+e2pRAEeyJvnOBfoLqic/OfLPor74hxgXubfv
PB706w8aKErCWADn2gs1CBsfLe6OVB0vtEJeYQiotcWyq3co4NS9/ErW9x82kWGA
fdtzECXAWJ/NuA/p+AST3y/stNdQI4SzykZAptwmKbEQ4FD1xRqoHwxQThj69dRh
7UiRpfpW7SgFl/jywtviT7Hvb8JKOIR3KLtC5R2F2SAoTMvdCXugvdo5XAci39oC
aat5gKi96S8tF7LLeyO8aRNZVgJm+ifPNh+54vxux6hFJvERH8fQfbiXHIVY6Vm5
uSwJb5iWLopNzaeDU0bSL9wuiiqOIlKLhKy0bZapu2x0Nre8rrPgatjScedGZPxJ
48ucZ+1TjWKck48Tfii7oy/EvGvLSnhT24g+Lughw1bDEs5g/bec4eRiH6A2iZzn
OCeVvXYDjSdQF5VId00oRRN/8V7YER3xSmnoHXaW1nbJv+9S0xzg0tTtPWae7PiU
UvPO9H/3TS0/stDgNTt1zrDuk3fCmhpA2OTF0oYqtLwcGLIXP5KEavM03e5XG/W0
0z9ovxcvcamKqJsuc9O61tnsb9SEjvFx5QjW8r/wMokUJO9e9t31160RXR80Mwyi
XCGo0jvsBuM8YQe1RSGwpxs7QkCJKk4pKGujfGajlyxkodJ5AeSvln1PCgPfbnu6
fNQ1KftCBLIAMzN5hoAeJu/1EY497ux7MJAUuVMal2R3MTb8XkCLP4NEv5LFfxaI
YxPmoARcvHrZF52ahEwIOH0aimJjQvN5/O7De6tHuVEvRhJshEtbaw8mqFCpOkwW
gyzw0+NtKbmrIDd/VhS6kOYHxia31b8T+381cj3ahRKMnxaN4V/iaSMpgVbUYjiJ
Aepz2p4wdKlDYWoDwxe1Oup7deBqIfOVBBmxff5imoDcks5qt7nzwEJScgdZyAtM
9l7J5W9qzvzZ/3YAn+pS5xsok1leCqzfK6K90uHoqunwDm8eUALmFxz3QooQd+j9
pBeShadGw0EaUPQj+OmukZ+aecJLrikNHbOG2ulqgqepUfn3o0H5rptKqwKtjVm0
jLHJL4ZlEsEJmIancGTMmDs01+WLHnGkLroVKt9/OVB7wkv+xyJyeBjn7KF3HGO/
0G3LElpF3BaJqS7Ccx0nq2CvEGx7yKLvJ0oqBxlzYV+sOtB0Di2Lcc3vCO6dkPLF
lAbMFcONdftVFesQfeGzvphyH8VDSLP74E2UkIPpCSXkG1qyoHXy4xLZXFcxBeYd
LWij+XjMx8DhBxHGP8mvsXWkO8jdXA7m5Yu1KbX8tvkSqPmAj2vhpZASnuniflmK
XdS5eZH7EdzLZCXnhgOWvh10zu7E45nEVurMtAVKt0EGDr8U5pYiY+BPbO5G84r2
lJ46adkzpa2Mfy2WABzhCJULTF1q6jeEcodeCa0mvDVCD6jQbs5+0NDWxp6s4VxI
sn2qCMTmk2y80lavmG+Ij8OX/K9LGFSifn0XJANoeJ+TSWaz/K8ybLPFm9Ks9YDD
eMETHZV+OymoTn4/Elz0uz1kWbGIyqBjsh2hVKckTfHZF/rle9PJjIfnZiS9UxX2
R5eBE6iSfUcXkTuyPU4YWtBi1hGPrV1d4AqAVdb7WEgJjKCEy0a/gSm9Qgo6sjBs
n2Cs2+GA2VHU4nUn8z8xyiEk0gd6RPonOPohxrSzeGLZvDXxmAIv8GnobqfNFyui
i+FmHbTfqf51NyJM0r4FDPc8R0GBTUASjEUmuFvM4qh0ntQp1v0pAqapVUUKifXA
3XrZs9hSnJjbWDcEG/K4nfNxZtNVR/7G5Y9IXucnDTUTOku1X2OZ7/oDWKyh0To+
rCH5VINQ1ILO4+IvyylDNa+qjLxHSFg+W5xxF0/z6uU/gHB/7P195va983mS6xV4
ZVkXkMOc8hCMbcDr/DbV64rV4ccGuc7s6TaZ8VCyr2lZjtctK8CFXucOsZmFg+ar
zpy7WGg1OpWBQ8S8LOpLDMQ+SpQ/8bsMuNpHkf2PeJew+djERl60OTRmK8IFpa7s
qmJ80UAxWfwlnDKmkJU4Cw1Vq5044/9pQLZydmkuwaW8HJ30WkmvTHw2mgIjkdn9
axKul4CdAzdKaARptWdmQ3ox8/3FcupEgPdFSaaxzCJaKGvNqZ9kRKLt251Y+Adj
TRoKOcrkydR3SMCXBU3l+S3VdGvgZlvz8/iCKFmZkF6Efa11OebhSIEhz7Q72VGj
LGW3pA2SlcvBXhpvShuaESSmc/E8cUoLqkBgd13E3e8nWLtzXmNQxg5glnjhVSHx
hp0HgM8jUUeHrOdiAsDKYPKo9rR9KAhopa1Ywb/uPHf7FWjSvFZdXTAYQK5bMkLF
NCS+RXnCARsZgngxx/mjDwUBAIDTGrhfV/AnKnUuzkMagxJ/8ES2otHml64HmkaL
rJARgib86xwIFQ89yFamYkK+/tU95kw7M2NETk8otpR95ilRIEeIvuae7bv/GG+r
VzY+3aG6OFXZCJ5i9pnIe9CKNvcSx17xmTY/cFpxIdoKN1dZEdEqlxDzmKHqeFyr
LBTJyZLjkj4NjDNqsQWRSL9CuA2zBUNaTixOq+nAYRj7EGTb+2U3msAwgUSabFmI
QCEuUuefcY6qzr43K0adSMJhE7h02nD0ryQpYasEGDCkWuvqnBWmP0hQqmcmUSy6
s2iPWjhL3GUqdDPEPJ8ku2RWc7epOizU1D5BEtSv278LyzR43j0AeT6KXAvTIeVY
S2vD3zQ1jYbCGmCMa5J+gsGj2Or1w2G8cu5No0OYJbQpy5jBtxoS0dcoF7G9fJhB
e8e0y0J5+uJL+RKBmnByvI0+TvKEMa7/DNsDRnFP2p0tZ6I9LtkgCpo5cQApWWtn
+cRAv0sman4CaUe2NaLCKHCf05eavxFl4F0bff2HGp8G/h2f52dH4ZQJ7GULNuop
tsyI82PATXa74ABkfe45UkkWpGeNnj1646GPh84TYxmbKFodgwAOTZSewSAnMQ1x
T6XAnu99C3785ArQ8TT7nTG4ZWAm97OtVCiW1LnQCBKCJcslw4/XFumaqaa5h0rO
9j3kzVahdPzdFPoj0k53gpcZoivKaXYOB4MmV6rg0XRZUe3D6v2JLw/Vl0BS4Abj
kkV//z77LRLWdRwoxaI6iE0C8wUl5XjdnkbBt9wtgeIyRn6hrJabe0X/C9uS0iIS
f7DiPKN5YZMFPde7jZmZiDGYY6N6Ym/VzBi/Xt36cRds0Uj9hwnKmeyayzGVPPqj
IQjWk72igC9RQg5MHDP/K2cQBiZfO0TTwsAK7YkP4A3RRj01p7BsthczV9NGhbtu
6eZls6dbFoQbepybmVcqV3u7d3a8erOTeCxvm+dNCAoYgNPTXwcBLG1DGdBZraSt
pRqwwvGjeKxIGRrOLvBbyYx56bipTw0xfwl/Z5ZTxNISWtJsT7V0fEY2G62acgRQ
Ca8xDS8j67PmdptGWvGnVvcpItNt+euvrf4WhHxZgC8MgTeMs0ppou5hNev7LFqA
FLvqNRbsEVF/lEg1jkFcdaLQCcoMeHAxQ5qLrUt4kzFJ481+R3zOcsAGMGRohS8S
VONRfKvsSTsUGRyJ1oXWAnQY+XPANIrDWAZZnqEJWb/kfVbBpuI7dQb7nL+Y32V8
zdVRjCD9CJwi6iKV3FKt5K6n5ZFsBvxBuJYsrPF4dvbEQSrbmI+GEzLe14lB2pgF
xC7xEuG0a0QKL1Kk07mgqkkq5rWhVNA9MAVj9qhwoVv8uJp1VCIHFqHnuFva0xlb
w5Y8YXxJj0QXauTNx/Vg1I7UyNpeUXlN0aDU7C74pohd0xmElHRAna/VrDpEMGjh
IKBNKF7OKxCSm9fbKAqpfoTM45RQPYAE9n+ACAEmYvzPttZp91hnuTAzUs9IDOGJ
3f5I3gd9dyI8ua4nqA0XyDM2h7tvaIwPOk3n9DsKsere/1LP7Lfd+79pHjmRTjUr
UJzTbLa15wn4OjIySa6vepjcnFxD6JzSN7d6mirhSQ/14+lWkgy3iSjBLIdXEmsa
NdFCsKMixkkvnnzzV6d9i8F1uWacs8HGn/3In6X1AjW78rbwPOfvCTaEALIFVdeD
jNZuZd6MV+zVh4yb0Ye2u2F3usSV/hNUZA5uIwx47gQ0QqlQ08v4wtEVWfz8Fbff
x8/yY6q+/4E5pLxokIrn4+a/GV0i6kzHNiYJMm0G+gOlBaXsxVJZrcKq19dfshR/
Yg+E1kC8qjr73HoGTvJ45wY74xUoWnjWCxvVEHsJfV1hTKQ8xy0M+30qTfJMAA/V
75AWbx8ZTdxzS4seLPzEZMYoVZtq/po2JprcU3vV4mFMCYEv0uCi4zwpRBbsaAVB
YXyORBc2L0Ke+lHmJRQd+VZqokGNec4tqEeUh5u7wRhbvAqVO1Erpns8YZztz3y0
aCPz2TYkR6jGbRF7O1x6Ch/66RrbpPT6VICsqqRDaIlqA7HB9YWa5pcQxJv8reaG
Vqhb20szmQWQ+d6fmzlMVDakOcw477LxW24Hvf2GN/tXiSzpQfxY1b24ls7+CBM+
AVubQdKdFXIreLWGElwfNZyn7xIkYVe9SYFBuZ/rtVENDSCxdOHfbdvw8IJYHdKG
QWpTuSXeA77MBlhYI95K+IxChl4c0RVGAaZPeHbzGBCmDnedpAf8mWnUOum+04lb
UU9pgQ7/VR0aIcLuLcuFEzkOZ9a074GNancXL08bdUJ4785CXPk13fSn9J2dOaSw
1bLIXPXCiwuHS4U1PS/scCzbf1UqFsWw3UN1vBrbRQM9nqIeZ0sP//ly+HOJqO7B
o2lv1DDgS48yobYZkkFahr/DeoTYPw4DP8mxcHZojB+u+8lmOnBx98ie6zCzOb2+
+oDmA2vJ+NiZbgwY1sDSMHK24wLq2FqU6qRuTusiLQrFX0ZtuAWimjc3bTrQUREP
dESK53t5Yr3W1XMRKXlw4on2X8s/UlaQBv26+EXhTJBVi7I5maNvxY8p+Hv+VvYH
MvRN+oFQhciWBFWWcoyaokDDYaRaZCu9dqwOLtOsC+rQWmXQ+i1XamvbLqq7pOn4
SN5B79RdPkWzqyE1n4Mf1jmc1U+k9zsx2QEZUq09dEtwBWGfDmufiLBkMT7Rs1mu
YQIKmgiNUB9hBceGFQw+I4Mq98c/NLxuYSGNMoNMODC71X85aEIvThT9tI4ct2kw
IuZPyKznKrVPlcbSgEpNWG0+jwkRZvjJu3i/228LOtiz7Ke1aMu2TcUkm8NEDCdX
/WzDStKZLgFdplgUCHTOj2R98Er/j33Ibs2VaKSJ3mLrxAY8ux0twan9GVGodusn
SIWPVibsd6Oc0yZZ9cioIYj1pVplBWnB9W7HkUAi0unMeZNV1vkYogkgv61ZWWEV
R3TUdhTSnfCZivO1ldg1WFqFEV21HgIEkjoznZfLqR4RjdZGr2eKzYVIu25D8Zlp
0N/O1zSRmGkR7GFsQr8GZ0HVsZoE1/65zyiH6SLGOfzmzny4ebmd0a8yXlAKH99y
VfdBaUuX0yO0Pi2b/+OELqX9/q3/QIC/vhr4C7LNU9UGXudc53OLRqamthG2csKW
rHzaDfbrF/gAVBsAg9UELB74850CaOm2ifmLoh3+LQTWfF87ZR6pTIG6igFX+5Ja
jcX1YrbR4sUS142c+bpCo7yJdFEIAM/DCiXR37JoOnggZeaS+v/wTa9kzE9AN6Dt
a9LgYNadEWsKRetZ2/T+HHVEHuTh+4GZJyTNlGheVjw3LnaNcJWHLGhfTBBaR48N
zLJy0yAjTqcGmaEup8m70rH9AJwFyJ1QUBDcyTRwXRDZLpMBCErhs0ry5t46RIJx
kfa8XfdhwXgeP+Y+1B3klkRoIOF7rJ2bJ6naO9bVq0884w5qj/AyS8xSxm+aGfcE
zxp2Fm8DY4t5eg+JgRWJxn0kh2aCNU57SzvqZ7IdT9PlscA0vN63lPwVVC1/kUza
FScWeGoYV1cDxz5lxyM0xZpswClU5Ta3mEc/c+qXaVOYxsHaakIXTrYE2vYPTAPv
4vUuz4gFHrweG0PE7frvLoe7zC2ZtVTz06+Djm0YXxbflJpsmAS3XRSqRnwYIUQ4
m2PbbP+1OCasdA9KDAq3xVXZH9GZawUTmHqmUO5HfRUUOE4z0VIk0YbHBFfNi067
m9ePcIvqX7669IeS5o9RzFyaA6TSVJXtcMq1PLb4iizBKA9vSGdL1VOpJ2kfnwXq
JTD+NYqPoso5E73xRY9njdMSYEO/6Mcdiot+gChILDE/c8iTd0c0+jsY5zhPhFAx
GKZm9aLkaXzVTbkC+xEUVAug4uXXbBN74kmq2pkp7FEH13ETEIW1seH1e1/j986T
SuB+IBWD86LIM7+FvGoU2pAYIJ2qZZlEupPQ2bbGoN57ir8ng36wKZPc726C+Pg0
36bGQsbOte9Ow/QTxwH6/ej2x7A25v6yrcRX4vcQLE3caEe/geMdk8tsCgIASnAK
aiONgO9+G1Mrh1rrqU6/TIhih6yrCBOEwsu2ILqZkGCwweRhOGhKwRbWkPFxNcre
2InqbaXfBiWKu/2gENd3gDOBTcAA+iN0pSd7wQmNwXYvtseqbFjHl3T+yQzwEzE8
c3jePVCZrJDIDGbJV9Uoh9mADGXF+qXxJHHD7R1D6Yv1K2kyFyi+KM6r5cblgWe1
fgFQZVe6emIngJmOXK/tluqsd3ZIjO0TMcyb+kuntUSjyOq/sYPei54+mwwgLrVe
S/jK5tdLt06H0/GEDmT8IjW9K0asvtNBSpACoSCoxv10K8gVQcxR+0JcaqT4Fdnj
erZeNau1RTVFMfNbpTyOzDFAjY+fQgQXfwkXLBtf56+9ndXHPbMlxaiLKNO8XWEJ
R9XaFYPMoemSPuGatKCeLPx1kWRIv17HIGD5WAQBqz9LGUrEMPax8LNSBqKI1zT7
hYocbQrfnDzPjZBRVQM3vteJcTwoaa9aSY0KmRqE2HfpILiNMQPxuvZwmNQy2/Ki
Jdvfe34LluB/9LLwKjdCJNe+iqRUWdXN6VLtydbzY6YjyXJSfLB++bO087KAb6iC
UCYgZIQRzaf9dHNQO4+aa0h4Zuv5YaZtx/Y+hCAsC+DoJB0sXt5PT9fxhE7Kg2hT
BC9ILwJEat58iQoPqcL2i8tIj6WyUuIf7zHA4PE6YEspD9Bpfvu5RA5MkvixF+z2
Ozsz8BHe+N0HnmfzG03ZDYBS6PPf7jBzzb3PVK2i5/SF+5ZASgPu+Dj4Pr5pSH4D
+imJjNiU5YNL0+cu0iKf9aBvUR3SvsPTXHIQ+lf7wpt7p4rbdJaO1MY9MKCVCJQa
YT0Ad06MAKqSSFTfXlv3oV1tiHn/+m+vn+jR0xh8PyS34bCu0RdqHwjqVr1AyC1t
I9AtlMaTwgLpTJSvVPbshvUlqn3R7KRjvISWILN8HdJ1+6Wn5zIMhq9QPSycbK66
XWqI6C9fDs3vyIYrtJgaSgCabc3VHZiHDmPFyOkHcix1Ott8JUwEFUFU+BFnLUBb
2geMpVo+gC1eiYK2xgOhBVX9mWr74j4d6vGsvBUSHETGe2UbOli/hGwHNBaJKlma
hb9idM8rQ1jb8HitoUaxvsiIZwMhFOYbEr8Dh8rMVJIwkGe9MteYgt9vp+oLIueb
lmLc4dvP3xUIp4qx4ca6YbTanAuWzAdA0CCSlEI7wvKv1A8NTyiTzzYepxIzHJeJ
1mX9XGbm818PkZbQFGVegw2PpoIuVlsJ0IYceuApU84GrNXCP4Y23LaVHXE/bhOT
8S8tS93CGobcdLi3+LIiUWP3WQ5n6jCZ1pfbtJWctVON/IqxoWzhfYxlfyYdd5UL
eQEgp/p5R/1RqcbacjwC8gx5QftCYpGPOB6OKuZvvZURo9okaRdcbLyyfv1bpCuK
f3srR/3rqztsjhu9qgTGjyHSZo46uXIKRoqgHPFMaEsMpi9qh2qXa4eu1NqRqAKB
RVGAzHc0NN3qdu7K59yDTkUMFGcQieI0sBv5TtCLWHBBHK9EFg+Od62BHsYA1bG6
lVK8JRoNO9Ve31ZxzgAVdc4rJB7cAoFlOJ4HFFFQe2cpsxR9Nb9ofkIy+gwuU11z
Ppi4TuA5xm82pTwe/t5esaAgDg14gkPB/yTmPthe/9FV7xg1adgLGIVY/eOZytLm
LFcT2FX23dYUYiCH+05ECBJjNO6ufAsOJ7dO2HizViyym69AT+zUeQWCMzodmxCX
0phUd08cj/Pn04lJoowidrjaajaFJhaXQ7jslnTx1n3mqYmdleceFDFaq5yxnEjD
/nJitZ6idqu6SooRY59KJsxymqDxwNKftd0sZduU7XdJAw6jE5wKnoYOqFOtyoAh
a2EVXxjUXSxdOvibNqmGtAc6sSPetwW3sW9JiJ3b5C0HvAJ77ImuANCCdO25YGkR
6B/Cap0earz4zFLcatHgCvl99jd6pzDIM8D3aw7NpN+aplAV10ieHHqoP3kxOuw2
+/nty3yZJq0AVKnRaBam2sFqoSRL2K4AEPFzDOt9E/toKzzGjBMPvo14lWxIZzXf
xhc/Eik3QQP9EBCvFPxPSMGtxkbKjFZK5vhT1pZO/5s6owFYPJ+xGoYlLxtzjQTg
q5OmCcHg49AVRnlf16vkezlHv5gvg+UXhHXm5fivAJt6WZFfuHEFGiTtZxoBCrNo
YJlitb82yCWXw6J2PKlDvDywd7Nz6RmOSlnZJC/uwwaEYwydcEk5bC6FtjfQT7M3
ON4y3L4wJQFit8YOYpWWfHbODHsNmiuVqYFTVfFBl62KpF9I/943aQFfpQ8feXPI
E7W19kf086ObNKsgKtEZUUTp8y4qOoWIYYVSAhsCXl7Msb9YGmnTj24G72pt3+Uz
3dCtfv7YyZLDq5xgxMUfVeFJ6mKoNaqZhnnaHcjBaLVW3KGF256xAenjKyOA45mV
+RDpNGSoLXbBYvCl+dYT4y7krSMpxFwrzoJdhFe8+xEgQueF8sofYiXhgFWctmfb
r4li6vhFUmLLA0WH3qROUp4iC/y5FTqot7H5Udqa8gbaXUtO3CTEn1OPKHriPCPg
+ZiCQzcUmhNOXJsWsGiuX//2j941DUPPmvseorF+/ZiKehv1K4IUHXLcmrs27MZG
flMU3TwhY1HFZiDPeDP+vbJTHrR8f7iDAoA5x6ieR5Mj2z9k6nx9FNAXl3dpyJml
U+IA2lZrJ+D/N06QYlNXUnra+I0g6sWX28JqdiXcjZgJAaqBY+qgy6REzb++YnBV
WcqLvDDiRh0sqoTqvF3RzKKBNhD24XTqyABw+jEPMVZI5Bwe3sSRu4bwBOTlBVK4
Oa3dWSQZCCiZDW+09AxhMx5XGI5FLzk6L4Ej2UFu0tAhj4IrrLyOL6X6/yWpVGYn
LPDyUqkKlsr/OwVQXheu5kfEEY6YTIbdWkoJ1wAxJYZrBAFsv4ngxO7JsH0wEzEl
1wHzVfwQlNiZzU4MeFxYM9zU1EbU3rByIRdVPVj9f4zWx2zQWTnh3axm9KuotC9Y
Hru6qYKWk1oHNyPFBkPSyHmjspSrLPQHA194Ran7eh9CTVBSehkqa+0hK0NARET0
Q3dmq4vmzt+jxP7glga4AuKHBy6t6U/V4VgeBJtGFVaBMptTwOJii0bbWbh4SiDb
P7wrm76IDt9137YtPrbFx/RuEOxivDViN1fI0ZPIhDXEgAeDiQ7uUtHuVo+/OdeI
cXp+48h7Gq/DHyXQscSRfkBYpPK49z5PgMdJ6shloK7y5oMKymCq+khfhVmiRq2h
FHa8Vp4UTgFsA0IClAdb6igY9G4CF+ovqg8nQk24I6x3G0iK2g8fqTZDleICZfC1
3YoLFg5gB6YxhpM47j2yMr8Tg/PwtjkeTsBRShTmDrmWETfaekJwc9qmkdbUT62x
P7u+DGSEa7GIMHsxApQSBwNOPhkfDdXEiT0rWsbFR6Y2oiI2gnZ4/azSTQfuoM8l
4nY5uucqlrZv8lRHlkzRAwZV1ziwbcRMDDlzETR4TmR4wy/vuqPzVWkM79D15yv8
4jfNsUlL0Kkqo/D9h4yt5FMqN7SMLnfzED9uzFyBM/Sh/LJCnl8sE3Xay2WijcDP
zIKl56T/1XDIf7sXV48tC5Qec1Alh2eM/IvrsWFNq5TCRFTFLAxvARIAc/FlqLfq
I39WnTwkom5M10XZtssSt61d3rvjz+HXuxuL6lWMwggGvRFF1FzLvLGueOUekzpE
aVzhAacPA4gT9jikwRQL1yeg4kyLRGv7+vxV37hIfq613UODIa3+HMYgHe/A2mQE
Eh+iCxMb4haqnXyTcno39VNHjct/L8P486p6qfOg80ZIfyyA3ujB0/Qr/nAQq/ZR
EyLkjyoXbCEPVS7wtuZRHoAheqkHB0sokjVFPJvjDFzUNHK8i3qPLF3cZ/NjG0Ak
JdIt1cWlFeBhJqaiAgPAkm8pRFIiB8pdxN70dezYTrBO8JBjikle/ryCOyn8NrIx
kTKlE3yjD1+sGr6hvI/+CUwDMU1DXaN73Q4ytZbH77cH6O3FUkUgH1ZDwwKEOjCy
UMIX9k3SfYIn38PhSHHoatOMEjqUj3JcCDcMnEo4s85MoOt7Qx0uUUvCq5Uu4HD4
VCf4esZPSnSmdrkdw/aUwgPitTvut0hq7pbE6K3tNS53W+9dBoWA1+V1/4ARqZTF
1R6YNqlEEIWb0Kr1GY05Bt0rJB/67OrpnqzxjC4NNi4vZLhD0zUTSZmyVFwFOQCV
SYQMPi+yCf4M2dBtXpnEp6R9jSFugVslHrGCoyWH36D4gxtJhczecmQvDpTCO3ER
dd3GjlARxQs7nZA3wqpC+LVi4CoDQ8VMlpxo3hYV4HcR/wn6LtfKfkLLXDI22naZ
A8xZdZuyLVpEoMNXHpzvoZcYGEtH4yRGNFA6qlWbgaH7Nm1Bs8Eh/YzJVChWOjnU
37eGg+s7O2Q/gbazbK09y8IjobQMjQV1CWPTZNhlHJ3Ag3v7Acjf0htX6xrvfIOB
xSNT/gk9v32BKBaCXbaPGe4+oUhK/xp6kXIfEu+nbpWlF56jyVKs3oHrRcEmMSi5
Wg9yUJfHsCLGBKadS4O17LGjhiNHE3fFB6ByKYEikac+yGziWn3SxQ4tom0kKwuv
Dg9TctDvuVabWq0RNJaMaSUMxrTuaTk+2kQVDnemTFjoe8Z34Iq8SDYreuqwLLQE
2kNSmg9y7LtGDvyBtF1P5IomjUbzIDuyL034tQ8rgKMov+NEFQt/NjG/GaFLcegY
R871b12MTr65lZRV6zem2R8NWZHDY2943836ZJ3SF89zwqzFIxYc6S/1Jz/b4jXr
+yH+kqXwYA/JlSGqDjvxVpvABEI2K0kUfdfhMkopWNm+dJwf/x41eDGo+G17OAyC
ChXRffGsVha1jUtkzaZ8nokOfe37G+AkddS/W+uuYWfShjUtXSFhBDPy7pdttVUB
8GRBzqwoyyFBbzLCM6bKXy5DzDjR/vMt4uPUh2YZdMM8b36y3g1cc74HW+pm4Bj6
4Zwh/xK85CjE/uGhbzqKoXGaaL9MbpmnPQPho7zqUp3L6hRphZltDPt/RyUagxuw
vxRn7PysQGpw97YzJjEIrmUtyGJNKNUgAwnDmQVWbo0BSH1QzPDoNO9WH7ON+1ag
8fRzw5IBJ/efKdCtq1cYguXgAuk8a4CyOMtPQ3ROtNO3mOeoTKPsUDbM8b4wMMZi
ibpLTK+Gv3ObnySat/xDySgrcG2/fst23KlYTi6mHOudmX00pj8aAs7iNfsoLdGm
FDs1k2BMj40GpQgGCphFj3UHRKj6zYXP6p1q3eONIzJckyOmE5oyU8eiW7CkwcQo
RkxPU6BAJOTruIj2iDI7yBd3QxUV+6P3Vz/WLbDrLamMqa/yJ3hUhPOfgLVi18yk
7d7DTMnTm1Nj7jlAgryagVRW/Ughbh0XkFqgc7wIQ/3sVJA1zM6+HyokaaOCKqso
7ZIcYp5GCZLeSoyzH61ceGclqGslyhL+U2zfNVwknbuD4kS135//l+Hcs35IhoEj
RNGmScxa/gj7QuNnh46YvSPPg4LfJnCbI6j1Cy5l6zMo4wO04Nm74JmdvjDqbTUw
9LAoskWXhxN9acbh7tdSQEHoh9NqjduVvbPJTd1PhUHUEk331ChSmRXopJdEgVS3
LssBGgAoBEilUF/3TjaoYbsG0eROrJlrzTwYR/OSP7tWzzRC64w9Byg6VjvNPjiQ
m1ZfsxxLww4/96as4KmljxzNcOpt9rVRf0N0bUgjTy8ANlfopqBuxC/vgzZ+D35e
di1HNFzBu+2RwpstV3VEGLvtCMlrdc7LHj8dPyZusqImowMms627udcUXoeRZjwU
fDBWa1s+JYMt9c5UiwePbf6D2l8Ib67pVyZI6MJ4s0fYiEh+bAnk+chqBCA1MEL+
HKqvZAs9ppbqC2EhRSaIDkoPm3MmKgZzufTZw1AEZRYzlTMD0zXvlHY2QemNgkOp
mKAk2exHdnNh8DKoGge3tqRjidu3DT9K+Jm5qyUGjp5fjmBHjkU3eYJ0jrRb3Qle
RrTub5oJ4kFtQF6OB2v4atk6xJ+bui1mXIW7CuG8nffjhTIyFjpbke5Kp1Dg8GBj
L2w8SE9SYPl/lonp+hFPwFB39xBzxNKnMGZ9IUxSPj2YM0a46NnBuTUBUFALrMtC
X2cVVhLFtzxlAgLKjPN3GiXj7nn4pnnEmaH9WMfDVpq78csZd8xhCvhoLlAQ+VSz
BeLwNkD+c1nWrtm/CzCUWwYyeAmCryUMyGV48lWGXWChCkfKDbG/VnLqjCp4Q1lC
S7FE5J3OTjyKAuZnKiSl4xNwm3uDJ9f4ZhkdJLEaQQYO5K/uAXV7VyW52IOfluWI
WIuGjz9+hrLh9Fmnl3ykyx+WnVW+2rPp8MRxwpgQspOtcMsdIFP7PEONUijJhl6o
GuSa2djV7HSuGwONpTFbrYUdlqATIZ5ScTBVVAKZUp9o6AhPqi1Zl8/Z9PMWDSzi
hJAIBcPKvYG5vgK2a8D3D05cW/bHtYoFBxIqEhddRh4M8KJYKDaEC/bMs6mgbmBf
gHENmzHVNkyzsl8TF2lAIczRHr7LooaMFk+HgAlelU8sEfWhIanJAN3FrKXBL3rp
5mCQajLuVcv79I//R4VNT64x5O1iCMLIMYwyPZqf2+fS6emfrAyHf/EzKHZmuL1t
UPhWlgxKt82dBGPfBmV7yOcXGrOzbw3nKB6TbuPZ/K3uMHFKDDL7wB2spV58KqUS
0oXP5buNwS+7jjuzecpe8VhkQwZ7QU9pFYKINwlxERv7a/GGksqXmFZV6gxJgpBs
ccgBbRj99t66RWEZjri7hC1Q7L/4XVt2OXEtU2PlN22sgiZw3Hd4Bypl2e9/2gfL
TaFKoZrzDbPcemVicykwYwn5sgprnkXhh9Fs70nUPS84VqMyQrIDjfZqAmxUIYbc
vw1O9DC1T2OUynclL7gGh+1X4eRaa8Dzg85OckoPxazfgBGpuPnYJdVBLn/YKG6Z
8++4D9f4/GIMQpH7/hBT72ePdHieo6gIA732H+pfB/jy6ANFOwRwYn+kkU5Ewg5C
uIkJGr4t1kl5D9NMnTGorLZUh8XTEuNBsvpGs14HAtHcEbkO4PAAuqyOmJQgGuff
pq0stDxNd8udb5u767u8DkwZkYfVnmVJ82MVbItKVNLVflZIg9kQA+K4cqRL0OJ4
pekVvWetfoh5pofEgZ4RXOUVDFYlHq673DJmhzW3wSWrC29qmGAkIyw28pjUe94a
Oiwq7xTZN7ui+QnnUVYv6sjGPbP1dlLMDm1e/riLPflYVaa6OR18vmOj5rNffpvG
Nl95t5M0b5NL8jjuG8RgEI1BguV71Vbvprz13ihgupNldW1tzULe/0qtTAHF8oMR
SXylYCdCT95wU3UXRIyvZzsGDaMQCww5nnPCnQ84hIUnv32LNkSUurBXuFmg6b0P
hsDZt6cuWxh+pcLznrhTqY6VzMSEGDP87eYg21wHNd5bmbg8DioKTG8H9GroqiG4
1NnjBogVwRgHO5xFOaz3CjdRTJCoak7NyXrO5hWTLSVCPG5vmZkrfi0buxlB0mD7
ypAmjHI0hhbhIPcx+DY6vwH7KMAE4bfciDKdpUfdjjHxrOhWfsUB1ZU7W70CthnH
bfhG/Go3iiqxdU28ZsyS12GgceVe/lRlxfDCOgIAuK7UY0qVuqr+VFC/QsJCIWS1
3i1aERh/YqlJNeOsn7CIsGbcnjphGdF2JaKJ1dwFnRoJpk50OlYcIXQ4C5ANsRHB
994THgDkZcLaF+9rmQLESGy9cBJ9ED4iEVUjTLOKGKZJ4nPIU/g/7SPTvPzwGril
zbv9TaDS3criqNWp+klhTRfJMqB2q6HcSa905NsMd64U5ropFLFaX/nvhFIBVwsB
81B2F+zoMIEaWb2IKMv9a+Pve/4GZuys96LM5xbUGshx0N/h6R/W4JgtPKHrb701
/9XpozoTPRDcGchTHFRE2NznXJOA3Ppd4PsF7zxVqYU0rwQg7spkT9y5DebgTVy6
nK9cavh2xjG4cLnY8efi6et1LpgOKXYZHTyhsAsDVMYrI61hdn93Ak4VmqYpCOAx
RkyyxtE87SaL7TBtZ7TZm08SSgniH5kiikslnUV9TF9glvvpzaF2BpC2gq+nd79n
TIdmhN/RO+a92ilZRTgqPtLmv3DSobBKLgjJAdbjb6qe0oiubXYUEEc3VNQibgJO
SvcpMDn+QoAg4F+uFQ2cHXU08GPQGx01Wqjer1h/uqvUsOLNR/JyTHCXRBqzjKzx
Eh5PvARr2nTsJxStc1jMuz5tr0x+9x8ll2OO0TF+H4Xhg55B4y9+7HmdlHfU/N67
HodSjUEiFWWVyzyOUkFruViiUhPyIn92JDR8oYzglLnocGa73/0NeKM/bfZIekab
p/eUPExo19btKFXMgNwn8299GS2Wwl4RNm/irrn0joKR3QMiGWLPX4nbTYb5ozgC
dVRe4kqEfW1JxhrrutQq9g9QPOby1Rpw3p65fLatODQUSHxlUd9SD578uMxP1ME3
YW9vRNOu29UsJKVUZFV4QLAeuqHEauIh6sIvB2DbV/lxXarOViRhlyF3jPlOnTrp
zN4mEPUCBJ4vqeR+DKv7nMz6k109S7RTghQ7dhfynLvhVd0Lciz4RXwUF5FDXiej
IlvS2gHoVN/1+Y9fqXkpN8KQMrEOiNAHD14Vcgs5XPr6uXWjL7VBevmVf9+Lsy5o
5mJOdLWxlEhWvdPVQ2q/NAt3VPQZ+9kVE2zighvdW27AWW821Y3vkTBBlxfkDdLA
KrhWt6j8G15tYo+wgfTbf25qw7UDtl+tpJvpgw91+PkBg7RmZUM14eHT7W1eggIm
St5Ees5q/OKibNSP6F4PLPkulzq9+REbxGafPv56YH2ZT3mR06+CP64lyu5mYpUj
2SNAIOXCw9Z7UmQTe8x6hF+W1sxVjAhOrCi1obR9LMpijeeSteHhuOQFw0ttY0d2
E7278x6aoJ8BeUdEpAANg9I+3Md5xi2yEArLzbCxZQzagsqTtzxO3m4/LOC4dXr2
RA2SCPgH0NOzXvcM+hEXzK/sd4Mi5eF6qckcpRl8oKMRMCJdejWxZ0C5H4On/JK+
wqdvK2P2zyfIcaM+XLkEPYNEu4xDt/m5YsattlCF9bZWmI6Bcsc6opf569ftI5nq
jsFcW8I/MphQuv0N7p2BwtUhjc9hgTsXEkz2qW+dskuPPeoJA3r64u/EW/H7kHj0
6re/YQ3U0qKsD8HfRoBRRIEIT34XuUSor2LQhjvJmjhYGUcq9lRJLSajoL5HDi4V
tGvf0NQNpxl2lFy4ecEhZ5I4F4PoriZed828E1s1jZOdupMhS1Cvd+XInp7vccG/
2DfOu+5tKiEAuJBZCS7EjBYV3bEc0QwxuMT9MIHJtj55YqoYmFqnLpI/ogfmppid
skHnN4YpniUnw88TvyKsU0vcaGOZJ43XeKVwNjvY3RMPSXjAa9KxFq63MxNPwExH
8SqPBvUPoYV6+3VQ1fHgIV8ZpOxHROItTvpTmLxubjxML6h28jfet9dFojsDQ+Md
Fg80wnI50RVYg09JHQ0/6OSimdfhuA3AGStfNbdG/bSbXIlhec2bgED/h/qAta32
4OFCoXiRngOU+fR8MRlOe48nIW6GQUXvyho9wNT6qHeaDo1+Eyt6s8CFh7R4hEEb
UdXrbR60S4Ry9fQu6lf7Wm/8IysSia92XKmXK2eUG2fTuUVe+DPcZ8AAjfbQLJjt
6T94WPK0FgupZmrWKJ8OBCDHBaSadbKKXc16Bnno+SQhPRnCYiC7lGdLfZos3Rji
0MeVxydSVPeThpudFL/uAYg8rMp5YIqgfIyDS4R0w+7OIDitNyQbxZQhGIpEOTKK
i7IK/xBQYK/mqo5dzHMTcXkzGblWCr0ZVeqIYl8n76yt46a/RgLFqrTeK9JBWRRC
XLXIHFSh9XA/qCMsJsU8awguKHrmTcQwI6ZqwkJXuqqfh7zfa2fNX2HUfnT2E0A6
JqbcDkXo0yYURTerju1IDZguz+hj+ys0ST4YAurjD7VQp+qT/PMim0PDWoafG/pz
84bZIGRASRVZ25SOYvz+xO+vppUk6rR8VThbyoLNjMJSACuAygKENCDQEk0SxRvx
nkWAP3iCfNoPNF9vGVEDgegHl249BVVh5xevilrUhmwqbu/eaHQU2EMZbTAi3cCm
9rdIqT7abPyhZoRSlQMxtKFkfswaZyGYJHjWrD4/zjfFR9tfr5LeCijGYW9wSfGV
UVpedkGfeGmimgdGjAOtLwOr4uFWbIy8865XtRIoUCi/jsfy5ZQxrTM3zS7R7MQY
Am5T6zBBuywzPF7xKd8wuRahIlq6ywRrdZKaUwfJC2nkwum9OmKd2wB6kWIfs9Lz
7PSNVoHiRJStOeACo92bdeSJ3pIfrld7vS5L0qSy3lM820EfWPahtlw56tLu/yaq
Tlj2hD/z3gmp+2p5yMU22GJffv9uxyhZn8+Rc3/x5HFYsqg0/8VNQiGE67k+JSIG
W7aodUsR/ubwDpuR8br2KVCuhHtmmKu67iLT3z4pqgkBp+yCsquAtJ4KR3SbIfDH
aAiJsnx2hR4j35DTnxXvpp3O10bq2bpAJ5KeyoxoZ1OQwpsKpjddv0OPXiKI6XP6
4db/PNzYLRpmNwWL546ZFvDL4SebPF1lRVTeqG7Buf5AkwWtYlv7PWU64e6g+wGU
xaLxY0mVSs19G5I4wiukDbD3w3lkQeBsmFq6yvHTNuh+htTFOBcVnXigsf2tPjZh
IuolKMNEU6MEyyAaZGSfQfdUgdcVHFNUgSFeIqAiRnu9fuBSniKueiCSSW9tzcgQ
TU/VAeCaky7SoikHr3NxU8ZCF/vT+6b7PG9gnLLuXoNSQ1Y4jeEP1EyetmP7z2oq
pLXquyvwNqYlKaj/vbj3YI+3f02HGPYmHMXwHNo4LB/z4WOLQ89ClUfIUPoFa6UX
x0RVvJF4wsexXbIuNeEc8jbh0UeYoYKaVgYTVL++w5dFijf3pBHJBukW+TktmWun
m6HYtYkJq0xjv9cBLwUSOiI+cTwCLCX9k+oaQ6yMfppsusjxYsaJwCEJCN5wmDjM
HxvH95+frY3y3fVm78BBRTL9Weku6hMIyvYShyKrX+GA6Plo/x/O6gqRYFUzsPfP
EyqL11/8hztZTkjnb123UMNiM4WeCug0htWt4BUYTPMJxq5IXOLHOTqWhFChO8wv
nGFV1coixH7JElCCVet0IPuNYbnbT5gp08CP0aFCOLt72EdQ4sWGE0g5MSrBz4gj
Z6rnM4wkR9a95Wf4Nx0UtWd+nfbVePkSkbabOK0XafQPdkDPgzZhpJqJ004Yffdn
ZUjFcoAF48Ng7wgxKmqhEVDxYyRsL7cmSsd0uRVIPIV4EsNUq3vjAhSt3R+XlXoW
I1KNH1XTiwOBasRnGL59bMZmMPW9fImRlwlN8A7GlV5owWIop0xf+xGHfGnECZy6
3+Lcgf+b5SsXRszBLrOSJnNvNyVTpmF8X7UrYIrJQb0sBPpnbfsJ2Euc9LrqJrPx
dursQMwm6f4jliZ6QzgtzpVEDeZ3r8BMLqq+I81VYdf+1thSljMupZFMVMascD+z
C8NmBUPbu+t2M0Ae5X9BJFjS+GiH/Tr6+wDq4yChtgpmlqJRocMyDSfSXVOOTstR
AnhEY9IBdyBeXLp2szgRYEka2aMw8jQCTptZeHbP7wyim+05TgkAcL+iJJ5Qgd3W
pggQKL0Jx6wjlQ54kxE2N5SLZyQAsy38TbHoeD1R+trrKwxhcxvcGuEfXziT89is
OF0BuyUIv6WJHmV709ocjQwF6uzi627DIouhcjCaaPg1Cr/RfndlD3d8E04ybp9l
i9EwE2Afx/p3wDgZpp44kLSNt2kB8hdqA5hJcWcw5zuukU5r0tjpYQD1HBbIiALJ
Fb25wyjxVoip4gZegpm1wwNmVtjVyaJW8Qqwn88YDavGD7WD+6HtIQIHt5ozOTCB
w+zSkMrdAsdSoTdMqhdgKXHkpwxqQb0FZk5PVA9R9xL9b6WkrbXUX9qR6srknryg
nHEdOXiEPDUfPaLeOlagCCTiVUPwlJllHoIZ1jqCfuIe1z9uLqxifL8X2LAptRLa
eRzTIKQs5Q3vcM5UfBdhWdjGUw5W81jGI2F/DbAjHcRS1ZoJ6e0hVydiu9kIeDVW
sH6V2OyGRxXkVY50pITSJ6qXJiJ2v9MUQVrFnWkWUySUPtyIAMLsqlzOFh/iZPOk
JNS8xMBTRLFKD4PEa8Gy7cj+mYREH/MwWCF0llxpEwPAQAHmm40vfs+LI6h70xLt
BHF27nCOWmvg1ox7LbsN7sCIrKRqQ0m19/SLEycoLKSJAfpRj9m2SK+W0EuDo6n1
72h5g8ul7jR57eGJyzuSVa5dxlJgkvPsU2F+yE8RFVpDQeyokmqEjvRxLOZahWhL
sqXrKfvyh1S+3/oqyLCXmUPF/vKmpU0Q5e2K84E0/NFJYkv9/F52Hm9KNpc7s4MP
dXNiCdHFtO0djSlBRdPxo6361HMWu7aFUoSztruZhx7UBxF2gFEhiBHTlZHF17+4
r8Z/RJsJCKhTSVDOCHPMecrv9WUPJPut7IVx2s1P5DIJmYEuPQw62Srjv+qdQN4A
ku0blhrsgq7Ag7nbTq5we4+5c1Gg83JgmeLDowMnwKXghWtU/EfyESKY2UebW2Zv
xhz4oftJW4IVDPppder8FAY/ohzAwFXThNFjxMiLLcgFPVgm9wtTlMMQi0MM+MY3
H7LIoa2LoJenq2PBIkoPqFgm//OhwjQRKHhkd8P9UCV5DnelHSSlSdC7w0zRlDc/
tUB/mYLDIeoIzP5pDikemOlqfi2mA9tV0mhiOrPacvEGr5ZSLa9hFVrM5epwnVEa
/z4+8bq9sOqEVBmBxRvQ5o47ioLGvE5FqMwFJLALEFi6TPAsOZBnmKGmCdBCOaaa
OkOOOYROOiKUXJpXlqXQv+Xslrjzgkbw79AAPHMALIFbOO1P5qTPV/G/i3lMWwNh
2KPrJiGU+qbM5kZ56p4oJ/Z5B95VE3yZqmjlDMI70vn5BkwtYs1V8SGrjFJvxeK6
0eCzcdPMy+f2Sky6HTEX9em/tDESTO4t0uvIzqDfffkpb/3kGm85slYoVzNH2Eeo
IltI6BZpsK2zZYW4DRFlSqTjZEPrwi09WhTX+1gGP5Za5fhtSoZtqvMMONtxEmMI
8ik0o9pQQ1K8OnQejhCnTvbHDfMbPKyVdSmTIMdauudIDarWwipIfB63x8jWguh6
yAkH6ycuyOiM/JYu6jKIRsFlUnMgCDIKsD6oPDftKMeJkF8uZLMcCz33ioOqKwJa
dJAOkyDjf28Ge0zPDQ1WJfqMC/LnR8QodTIPvbhhhkPHH4+keArRawIP/63IPwov
nU0oJFIAMiXmUk12JvmzneekKRmS7ZrgNAdL1gHkoXkGF6O3Fviqf0za3P3z8Z2V
9+N1l+HD4KRP+umI9FtOXs5HYRMVyXSitdceFeX7lNu9T8t13iJL7GbZdw0ftBBw
rKdNPaEmj2VZ4YxHtfxEdGEpyjEW2rjDQ9539ArcnJwyVqjpFu1m2q7C92NAluKE
1phdjibQa/qNiagwvOcLMI3tbSc5TpwA9BPAPJAFoEvOMcSS9oHZLffsFXAd9CJu
LLPps9YPFonRbcLb0t8rokC5YMgfcE+wQ/HFN4zFgx9Hic3c28HIVgyIZKGhXq1s
n6GMMUtHOpBfRH/C7vchC2bNEq36Obaz9c0F5BwQbyuRNQZ1GrATbkhrbO5Q2a5W
Nf5GNY/q7eXuA0LF+ukZxbusNyzGh2O02Qs58EvNAvIQS6b6bTn7jkQWrVz2UMZw
Pb5DofoE1ddbfNHQXt5ZOCzQcLIpkdPyEj+933RVmsG9MFQd+N1sAmK+yyiqv/1Q
AI42IFjX6iz7zAksY9LKKV7VmwwR0iHtbGalTAvq5BFWUUFR/TvsB9uc7EAp2DgL
TicTUigTEuWbaxkKm4/F1cghXHZZTldp4R3AOEfI8hnnRhd5xFLoudwmsyjA/QGj
qhyWA7FXfuobg3XECL0m06FuYYohtBLpwXuMXcZu2s5EuB2K/Hgi2EQnMJMLeMmw
KkWh5/O1e84SLK6/lKBMAJrBx0KzxgGo0ArL3hqRhTuw+DdWxufrsOl3S7yqDpSB
OjXbKDv8cgpyD2/YL0zfTQvBS9FZy+2NJCCamUw4T00W6MoOTndB8x2pYcytMXcy
kLZTHu9bh0gyHHoD7+q5+Wpasw8NprZPGrimsFIDbeKQu/mxrfiJ/ae4zo3AZvNy
Vllmqf6V6hMGUFwOrnDPZ627FpyOA+kovdLcfXqDteQa6K0i2rKqUyggrFkwa9YG
/6aSddRzAsabcS+dhM1IQ7xSGZylhfy/OxpaGkMqQdNDwTHbAlspMwTxWmw5PHCr
9WH48wSA8YSA6dVkfnNvnp6n7sErMKAHB07pX1/ElSYMB6BfGVqkhaxV/bI9B/CP
TCBqp7pdIBVB+bFQrlcAHgAOEs3ZjcSu0Nc0XmC8MJHoMQpvJj3aeKMbrNmzNW4V
60nJSkEBzS7mhYmsfULDx5WVDSUzNCaacCusMTV1vvzrnP3VcmdpL6I/SFqSGZLw
nJeBbgl2V4kxZSajKFELEYmiQFZQZuHyJ5y79WTo4D+/8I7WgTcwCHeCkrwmxFtM
/JRoxJau9VmnbJlYdTTVLRnsrWSP2d0IonqHgZ08d/Wt8nBamTlciceSvy4fLCAH
yIbCt1bv9TVaGLUyg3fTXgYdVOlH2QQobkY0/FV5C0IxVo664EsGFROepj+HC/WI
874mDDfl2Qgx195VTjJt7c645tdQxB4DRFa8qT4puvHz2mQVtJLf3OkDHFrdFtrb
11DS8ZiM/TkVuqrHRHafTpVjcowe4YJ/NamNx6VM3g6CvUABJQYQ3YapT074KP1m
oU38PXCGu+3togTWZiEt37YrZ0ghGrxX2z6sbVjRBt9aFhjBXpL9iFQNQjJHBe6q
nO67Aye+NubJg2qGzMapl4fQk6d+dFHg5Fk8AfsdECo4stywWButoqQCG3ukTdQc
zkRhFmDTtPSAH2j/gz817Jgel3igIp7KC0RMlgwPXReQLvh+ghmbHo6Ip/fG5nhx
0q1Pb3W0lXmhoyUL9ciLgEZ/ziMkCiaNJTd51T+YVa3+AVORSkd10vHGJPEgnVGC
D/o279a0z2cRrkWrwQrHQ+6G1ZHUM8fMk6tBVbowTfQQwaI2H1s5HvV/Io4/4v4f
K1+nEjtOjFZ68yLsLsAzBthxQJpkH7TF4WhP/fl6lAaDLF92dsd3ooIN2TTUFh3i
hUgHNbBpXr5WK40MJpkZsKbyBgOdV+fHGBpxl5RLLhNjVUG/imaKSFnIiDDXvuk3
fJzu7i/x98RArARTY3NQJ1qh0xb0UHl9Th05D+WzFH7hiER6au0cMyHwi+wYqIuQ
PQX+AWHBOYbAzQ8Kzv02GY8yF0+BJ6HBpzwlDO6+1DgIsZISCCL3sL+Guo9hqSJA
ol2FxZ0EgtB3EV/hRtp8GqwTHp0BjB7u2yVz3Zpx2s/8yeWUti7QXLiVLXvQqKvV
7IptMBWPslbVdrcM51L1BlTj2RtADp966E2JPyZ2vhl2KuCRFuFa9ZJ7hUJ5qes6
Uqr2CvBJ8PbSNAPTxX2qXgfzaRsPrr0WzShHuSPszHyn91GcBJwlmCDFKl/AWCUJ
8JNRFyTOUSPlPY32z6/ffcpWwdv7vVa+/IB4C8/MMLSubW8PGkX/0MhxWImhhWHo
LrsCL/8LCBgTwoOoEBX5fXdwPi/bgwaoNJJ0wbtaMeEpBvSl5ek3aglSZw8zDm/W
XRRvFTk07nI9IxC5GxVIDJBKWszkCYmQ9N5s7X75bWmDhrKZGwPxesMLrcFgGqrG
b92yNhNw8j+a4o96x7+saGuPfo8Jfr05hfMK0tE+SDb+Tcs+EdIriENpj4DTq4w9
EcC+mtW9YgT7gTYxmXCRFn+fVOryKYu5QPXiso7GQfGB6zPMex9mg5stbaxiWSO2
UhMauw+r6oT8qd3RstKR9iVnVjzs/JP7HV1zdXHQRRwbnT1gFb7AgnBJ4IlM8vO1
Lro9DZwnGPNR+Y904r2b5iileg0k/nU7JnDLe8lbKhUWWVi4v0JV1X+3Mdwh44U2
Rq7Y85ymtLqn7pn4KfIn9j4TdsE4/wUHY57NICisuaS0I4STn+aclOrTPDZX06XI
kpILb/aCHWLzFRVhtlgLF68Bt13vZAoh6Y0OrjbThA6viiCo6n9dw5cebpnDxBvg
0BNtft3j1IkPuU05rFhAT7C5nEy//AnQolhqMU/nPLPa8OhnWS/DEKFvcRu6xljF
SYCOPcM9ry0JV22MBK5IRfv8MHPayAw01U5oY8IuO08OhwhLfLGw8Qy5+JNpHzt/
hxC+hWPrvpdI1hNnjFOQv7DDrSIRVbUe2EmNmVRmtMSec1ypTJVcf0A2LTL2fIku
zKe+iMCZudDCElDLplNHAKTlLeiX+K8Icz6BILi6Cm1U6ar6nLmzAKRHS99vFVdg
J7s6wliD02U9DAhIB8n1leayP799lnX5wNybzPh6hjLcbh1BUYQsYOvooXRmGp+E
PPm/Jir1O+AsJn/Jr/wsJV9Llmqp5Oq0gY7YkpL32TZ7gwDjFBSAx81fj9I+WZcV
IF8eG4tJQ/I53BRi6iFEj3UqPGrINsCRWVWwHY1tykJ/Q4VnKfc1Z1XpOwAl11Wu
wyBeJroriNWhHMcM0dV+2xB1ZYF85ayVr+N3gpmahTyiH3d9ErV+Kljw4RxhQdTG
3jNUo2A7STf75ZhnxFFPzkDQdhoxBwRPC1/HpKSK+unjB1BGc2Df2LpcLZfFVVJe
PFCXqiZG8XbAz+mDlyx7jcfpD+SfxW0k/EG32aub95UBXO2FwJbDkz2GfnAY248i
7wgJfg9w/n0/B2zJqGkoiiJYNKale9Nx49yJD7p615r2VT4rj8V+U9cL6twlWowd
VJliTc1Zo8DCvAytwpQTbXg60X3672fnhJTh7Dsw2TR26aNMrLKu+Il5OOVUnq+6
iou1wZyTPXvkHC7Iv8ak1cxNLcZkeNPUEeF0klaQZCnl7tDA9+4YN3evhYF4FAYj
++LSGzGWjhgaIYzGvf7lmYpMhO3j70GWQoLokxn3fLDCy0jke2tixNFaSO2rnuNp
HUpIXFpqVAtA2vONtcDS9umIi61aO5T+alMiWWXBktb3+bNzN3xIaph6IG6cJ436
7B5NTrL1nqiL3iEvQCFrU0gND5Teuq7HDsl0jPB6rNBYCx46geb4HU9ZttHfGD+K
fypxWPG2TUZnnZRHUeyLdNih06O6f44EkgKcg/L4lKbnvx0urgQYTl2ZRBYEPhV0
BNnsYF2RrrtNGkKYfm1GAMtHuwiTGo0WaoNyRp6CoO3dH0kFR3BnNPJSPdmTiR3N
t3PMumzmyRqt55/Nmd937Vszcc08uk0ijwtEn6IIZb2EmrEWoPUv5C7+Jy8Fy8GF
LZ1+tt5Kt3KwigbFW1L1l8XVY+B4wtMvwoIAI/x6ac3mi8jEplh/MQgcBprApbRA
8i5cW3h1zTq3uKA87VRzWRxAtN6zmL6ZHYxusfUjJBxjlZkQgUDrqVWtNp5UQDSl
3uJqpqb6e5ETNUolznrYjZb/sjHKOPJD7X3/fkES9DoaIGHvS53Ia59KPyWmIRpK
SEy0DybIvBP9k1gNxt9wtvujKIwaITrOtea6CIttZLmfCQrlUzTeGERSn4SZFOKZ
oWlZGN4LTAgZFXQJWz0WRhpvR+ViWws64pI70yyHxnnHf52Z77cW3C+y7REJiC9Y
0TwGN/D1ioXX/Lx5jGSB5NsWlnnAe6umKmoZFykGs4lw4FzmLIFn0rBuBiz/CA2L
EwhwMQtvIwvIqRV0OKQy4kt7jJsqMPu2fdnMF9vZhwPakA7FomE/Yg9seeYrDqfv
Weloe98R22jDyncz3jEsVfD0bANGSda/UZxhUSfZYQgHDj5v94e67aaOIlwGuRJS
oKVQBXMoGQZe0Gn2bF+N0zHEI/JW3RyN3tpR1skAzYmKSZePiu2hw3BpX+Rm+pje
Pscvse7oijF9/27RsfnniQR1Qi8gj93wYA4oaDbf/qZL8/EcBImSVFwzvk5AVpE6
bKprfa5mK2qjN/91HrEMDVUNIXJ0Vi3V5nP/dWekO7heqBw+kskS6y+hyCqKttu2
piDaGyE7OBoP0gO4WxgWll5PfhZjh+fG6DMg/e59BqkfXOV6BcRAugBfUxI0zpO/
BuoZGOGTZSJCTmEpGatsQ3UOW7qrvcv2EOpkI84U9C71/KeyYmAYo77YIZoS0qIw
Aypqrz4fVNOn2RSDWNB6gUXYE6p6DHLhPrk6/ZL8ZNYuBjmu/Sdh32RdabyBIsJM
25I+9tKVbl8IF4hNwT1FhrdZRd55qa1jfG0q3I/HtvFGMZrU4Y1RcuFjvP8hXAl2
5X1Hd8w3KWFAAUmvnidJTf1Cxgo+bLM987KNy40o/U8fEPD0cLiM0SByT6fVLo3s
A4fZHnhZIROR8TM/JGAm5ba51ZP/0UvqWwemccKbM8M3FuVe/9ZR4qzNVFU/SaX8
GPMDqWW9c54vjvY2HUcqdzCwX+j/KBLLQwW05jrldKE+pt/RfN6ouMxh9fAPGpfS
ACXBE1IQ5XnLJ/ZLshzIsl8JB3S7t7QN3bzfigOHrFfUM/jS8db7WHhqxsBDdUFu
ZmN9deAmTorHInHHcvc62nSu5zQAut1wQJmX6HLOvQZq338DS0cn2rHbZLi8z5ns
nXMHu+M34tsW8yFsv3s0znFjL8tnU8PoMVW9Y1tK+tcgKCAZZ3eVB/9i8fmY9LVC
ykLbHkn117tLHx2hsf39nTGbyZBtczgKywfHjnOpYil3qdGiPoW1YchkdiAfU1sA
3iPh2xL7IXG4nY3B3Wmmtsjxw0nKJkP7yZqZ8VJdeFzC+0JiGrqU19LFdNW8sF7Z
XfpD90Vv6MLFt+uQFheqzT0RfppqFdENPvz8gvmMoRMb7eX/ZC/gYKW/S4pJHrGb
9uWUNtsqvdpDVyfD1R50HUJfsCIpOyc5obr0N5fIhBby0h0ZUrJq3pjKcLdGm6X6
I1aTfmqkdw5W+JeH8LfeVMLOSq41Ta5Q3n50iKSJf3wABpN/cnW4g30MJvCIa5m/
S2veAW/6O6QgH2xDsSKJm3k9K2gMgfCwgXNV3OBu9VIGgco+g81ldP47aEzBsAfZ
DWEp2owhCA6cQRkmUePQ+tTsCqAExsAwDDUSa0GIog9TnZdgegiiR+rGvt14J+UJ
bVOFDocY9FzXgWrSQn4blaY0p3lQ44WR6b+V3vKrRAr2dNLezWCUszDcqqaHLIk2
FRyG3Z/5zQuHYImv1ojWZSz6vXU8wx768UanKHL9WP5iRDiq4tCqz7N28a37fiuH
N2C5xnH+yjYOPyI4KyHfRhA+VxJaR2n9gpL6Tn4ftJxDz7gn+g/OHdTKpKeKEraF
Jyn8L5qSrmx6kuM5MICVjxWXN9CJazM71dLrsUpSaSQ8OSBwKa/EwBVCTm+JNmZK
aVK7pdQ8bG+LjrdbIiIyjBy6lVzEmuMYF1qFiKzyriKK3EUt4J0Hj2gBsaovJKgH
LcSVe0xg1mMojmBYeYd1mq3wKGuxV8nhqUdhIxHcWkih3KH7cD5Je/xZtY6WTcYo
SzWWiGQ3meuL1RiJIm3+epEzvfDWnF8cHa4rJwSA55wp2DoVYOi685bms9z3wb+/
muVO4kb7acnQ0OpuBLTgLk/8tTY6ik1/kW+MW2D73uoBNGslH11xQjnAcsWA+7Wj
1NBWJa3qHsTinqkZRLVGFZeCCZi60Xmw+K3ZMsUkOcXmMu7B/QWxoX1SC2EFLtML
Y8H+iL1CIpkSzwBMWiirhwWQB/SzVAUmeLanzTp2ZvFpq/O3ByeMIt3vaOD83+XR
VcWhjjGzkkQ0DMq1ksENikUZXDvdvyq2/A47H9MSYYagIMbd/BjGch0yGSDJbC1x
1zpzClhmCdhNN3ItmlVG3TMlFZroJQb/m+R7TIfWzO/K2LOS/1C7frQ3ztKX/L+R
/BBznd4Y7bfhC5cUEBUyxO8rk0hum9az2tDZjmT/2T42ap50f8wCszMBhZmxAwaS
TvWHWrR1ezs0ru9X4OwsrePg1WhnhkKyfA9y0QoaFZ3Th1dtTLh+lgHa8BBSXLGi
Hp2JBHg0o+V1fuCo8MT3C7yo37AZUB8ETvQJBMvqwvYZoexsfQQfBkDdMH1QovYm
7jlMvIdYYxhK+2ZA4OEvY1PRaK3CEoMPvsFdV3VtzkZUZAGLzti+7X8LXr6mrmmP
DJ8U111CzLLWllSpOUuRg5ztbzD/PU5f3RNpKpHDxq4E8iYr1DpPWarFLv8DGzLD
6kfXw5L34UITZkIUYaQu2w2EEgJ7pz9d4slFCLlk/B5+FXXRk5msCvdDHN4aQr9U
YZqgRDd37yDli1NLEjL+g5tzsEFKh9Obh5Ns7eUTtzMdKn9sepSoI5qU+zrvNT66
OM6xN8PobcNqD6CQWH4Z9i8xDh2xtWHkNliDXvxb2nHStNvfYBNa8HgQWzV4FSuy
a3wjoLx/+yjSgBPe7w1xrz6ZZXqpsNBVWA3wGaw+D2dz9GqJIWoy+UITkxi+PyCW
bCJ73yFPVnPa6pC/mg8AaH86xRPmFdw6JjmRUajQtay895DZ867Elyd9DdIyXXNy
kSqIsQrvRjBwF11JSp5gY52pv5uQ/4wv1/he2L7fR+Q9AlBLOVYzUqHXJ0pJ60G1
JJTwLjNbbV35Kb8lUvJvGJFZozynJunHTuzX6S9Y6iK2CFOvnmY0Xkz074sSzXAh
zeuSou299gpTNGQoxSh4pWPwnmj2LVHL+Xv5K+hICT16dIESpJ+rz5sPhPfqag0k
8xTeJl8P7Aj6YyJyu/rSh7RwwOwjpPyyIute7zX5u1gHrF9vBWfaQu6xW+z7sliJ
aShKHcb1sk8R6PrDqacHfdRYG4jJ8X66OiEoKEzG6PP5JPVUlWrNss8u6oiSPnug
Ds/yinU6wex3jU6K62dYG87nEf9ogG4IaGhIxacA8a3UQQXVNBS7hkQFvA3RBOCq
sMg+7RQI5rTBy112Eow1RbtzO6VruLin5YB5qdtnqD946Nl0nN3ofx+glb7Sni24
wH0/5mBCXbnu+r+9N1RA5GYpssOAvaWDY7QVo5uwKCfRkZ+DnoiKwPQKNZb6PSVp
pBVgZhWPKMJg1iiqr/AMJwFBirZAqELWW0pcBfHWDXJEhoQmE9nilfg4sNIjAc33
2XLf0meoYyQFuwpDJYAku9KisGTG89Z2B+9BX2sgA1y9BhGogYWxu81AmaovukV5
FeS8SoHfAQ77dzGU6pY/VuO5ENY9VaImvYVGuu3hMTemMd8YdxyaD7E9YcNXOWWH
mz+OpzWg8Fp9vMHlp8b9rb+F/OamsJ7UhGpOj//ZxenGdMkR1BOmIh6BzmAJuprE
2r/afdyVm0ZWoFis+a6NXL//m4Zbh30YkQ/GNjcA6THan9DzNwucFl9YJu11nLuu
RtsX6D9NHx5jCMwnoSRsGqiPC7VXaNnyC5/YwuEjfLVDLB7e/kjFy7ETaZOgml8Y
1dpNGtDPZPVrzrXeq8BDdYkZskuWUxIsfViLQA7QL+7jqAnBBjm863EkD4xElLVC
IaqRQEiPh5RkJg4Bu1XSCOftJHva0rYwbm5BeR8BQiGwtdySGUmQmwlqN1iJYEHN
IgO1WB/DdwyME5J92frxq/hrzGMNR4z8WUIOUCqVKE8qFT/9mnNrPPFgRzV0mSnm
cIcJEYQsUn9L7QsjSaQytG9G337UnGRgpeQuvD/S8Y/XISicPINntYebdc53N2w9
T+7KdoR7TzOIa4b2fbVA7tMiKxYHOtRO3FCYCWn6/4HkmzTBtyIprpJQSTDd+/a6
L+srTd8K3H3iUxaHxqav9ZEKCBYEfGtrzNnBGdTO1SADWBGJsT+IaJ81u9wzZevC
amLuL0zMhS/4wIKBEEH8o6XeLuQQUwesPC5B6d7Aq/PgYo1JmOofriwD/ew1z2Pb
wbzi6u5p9mKcwqnXEMZVe/XyfHu0kGipzAtELJsYZcjMjawUwpzRMv3wev8wFqyp
qQSuB7SwQK76YKLIJFOEwkqTWdFVdqrxtuHKdKnaZSNHcZ0Io4i+LDatuOYTSYYJ
moyxbC3sBWIqmXJBHCgO6TKwA+DueE/8c++or1s5H/8HOt7nWWXqGK1vyzVl6ZdH
L9g2zTpdqV9zbkgNxzKx1N/Zc+N7g0zSwM0eJPHBCFMI0TuYLbTkVRAFcgyRYKgZ
mVu9enASmC1D8Tu/xnM4/GQNIZMGU7Fk4hQvcB4A2BR8vn/nifUXLtYiuAZIJfFg
WwceLXo5CvdFza3tYcfz7mq/XyhePM7HxsFBuwHVzzojpmUbh+h7VOgNWfqCgy9Q
gxzonpKtXfOaD8kSwhuDWrkLXhB2rnPhmHKNWTZ1e/9zAMAl4pauaK60y/TcR9RF
kBkZPyPkqrz8TBGx+mO6Pa2A03wp2IUmGWUmGFjiHkvEwWLxxuoMEDATT7B15vYF
viCTjJSJrc4RSlXMcAlZPx6qJ8t/OY86z/vSrLkzBVulS+rmdZ5tGcgOuMGJPtD2
2F4EDq7ztFoCnBt/aWoT87HdVs4R3mFxS9Q9J6KNBuGGoZcgT/4Y1nx8wDDMuCu+
AZZgWmWd72NLfWwU/hvPEUdpMLQ8u1w3I6kOtOLT8HDOSLh4N6sOWqP+nyYBZUx2
QKZudt30kLS4yQ/MMvLVckeotlyQ0MZYToMUx7S5Um01A5/9DmPnmbpjFchBO/Gm
SOZCz3ZCIk1nAfGmEHm1siqqkTeMeyz1cJGCwrpPnIbycCnSvNpZznDVS4qKeLq/
mjXDl2nfI3LQmVa3WG2hLlC/4JwPSZFcjYx+iIhhVpBoxR8wCnzTl03cCNcmOuUs
xCKPgr9GxMmBoAl5ef5NMFSYH1CAGDfJha3WJ3055dlJQ5O35sI/GtpCKmgaOjIo
9yOwOj9NsZsnwxHN1jLRk44Btc3Pd0dTWZ0KU4KyUDDP7E6BlQW4ufr7chCmmrML
2fiGYWn8TjBt2GcSr0WIEvwqY3U6rOBBtzxFRanfRxOhKYKhERBdocrSe8LEZolP
UPJBch6PgLYr2brM/qTYT7OLh5wKlN0CSLa9t4rfbut6zVUMMSgq9mAB2uykcDnZ
henMpVbNP1VdsFk4bPYH1nB4NhtPX6EJNjT1W81teskyI/0iMdMZucAW0at/rQlM
G/OgT6iO895u5DIeW9O5Z1tmGzb+RFIuJiyzKUg8m2NpurTBsfEQrDVHYsKPr5Ei
g5flroXfmO6DqkqFsRRjmBOsIGFRlSGH0EyFrAr5W8vpgKLN3ylMTZ0k6h4dZ3zv
1jzE9lEHuuxcFt10m1liZqGZPeyrD1U87qzgIVZAr9XGs+ZPbqSY+spC4+b31tui
f0wYzbYl3EMkSd0igUXAyeZ5eU19Vzx4XAVaDP8P9hK3gkioTQlSBDFtlzvkO0S6
j8rIAa7rYygTNutx55Bvo/BHVqp1woMPtHUKG00iVC0mSiSjC0YEmJC4HZqU+y/y
8hTeH4e1zIMunJkFh19WnudrDkUbMtxMuvXww2cHuCQigQjnY/mkOaGOE+xfKlTJ
BZyVtrF66h+A8Ki9XAwC18gJXss54QVXX8+gbE6HvgeIn4siG3CvCnM0ElyxIklM
1OXM19Q7lKiueSnDiJhTfpFc2fLDpWeL4uxZIsaRuK+XAHoBDIj/cuXA7YPfJ86g
KmyzlRPl2XG8Zmhu31m7UvjfM5HzDHtr8WxgAjEfP6PqzMfKhIPF5W/CNmLZZIUz
0gNxRHNvP8pkgsLft+kFnNX1oEnMtgfK9C8EeAOTpdFCDHtW9AWJQmz/obKPOoEC
g4u6ehoynj7yizzQlmWn18o+0Xj1SeOxFb+N0XtRkyizvhCZ+5LdaTlPy7QE5puV
0pFQIPQLXWnZ9JavobYawSQkW3bBtyCdk0POhD3K8he5yqPKdfLDvH4gtujLeQUc
vGcQ10/EGhCBlGusuBDrElt6Cwg+aH+InJuoeg6YOXvrRCSYo45PagBOcTTmrMyg
HLk0wFxNuowrzpa8yyRuZtzsoZ9+863gNASYRbJwUSQTZbanG/HtAlEnVN4rlCEw
S3nlxI6iddrWUdTnpr7scz3LJ63EZqsnxRRQcjI+ajsjO7R1MebLxs0Xgbr0KOev
xgsGEEdBEBkEbHbWW0CjCYVjgSVjO0VxignnDxfmsLAnN7+TJXXAr6OBlLxlp9t5
dtBDmPX3ttyVnWe7zD5IfA77yx6THGvtrG5SOZ4DQZ93rbiPHIUCfxXq34aFXpym
lkYVxIbgeiA/7v255oPQZ47b2iwinMoygNwFGh0GRVWcKKJFT/PCV+f34ckCikZp
74XsC7Q82Ut5bEQOp5wGUgolOdMGi9+/qxmcLBEPVVY9wnuviAJZau6ZdOprPGsp
U/3tgmyJhhKNx14LO0OX1pZuO3RpHhmxS8QNVc3ykB2/RV3O8SQW3/FLVS1HSEww
/enUrJcusi86+8FUGfAipR6tWOc8Awrts2SbvB0L2DWgwYeFoS0Q6imdf5fMO1U5
XGFzK/YuWw4NxU8piNivmE04BxDcW7qRZhvw/zmYXe19nlIQKZsF6j8GUOqRkER6
5sR1TJz9OBaZrDnp8WE7JYMWEUTGNZqkjMER9vqOfcNEHchEMWgeOUkhthif/9SR
eVxfu6SjAxr6rnN4xoY+rMAQG7zUFDEBkGmj5nQf315rIKsucc43RojsEyvNJylp
2Yt0j1CAY1uWkNGibVG/j3zfUpwjczgzgBPjXJBK1exijIcQw8PRh8A2Mwotwmk8
TtP69EYIujowCCdt3nPjQ7wGba8xwHNonSZch8duL6JBvYKOosF4nffqq+54tn59
ZVPPYfFs17NNFYuodZbgr9dZnIBq1UFxij00s9DZzaCg6RLU9Faekvk8xbNogXBe
p8+zEvbW4gLVb2LRnc8h4+/p3H/p76XwAdmODlY+MncZd8BOaIOwMtM2169UQr+Z
NeBSYjNoaLrndEw5hTze4Q0jQEkyo0SCrxOExLAce8TNdaDKOaPAnXOOhw/C4ReE
2bC1+FqKnfbplRMJ7bPYaDXe3IMYFrlLt039TMFXSLwSISrqs2mR8GF+zgAnnM0t
StRCNT9RHR0M1mAq9QDBvMqW74w37Uk1r2k7fNgVCgLMw9terVI8TfRwpApvMaiw
lA0qv0FxgDV/l22+vnHq1xDyCpXWcdbiPpyJE6ll94wLcoX+NN3sLHVKJ6RzwWVa
DlPQoFnOyNaJrXWa+SIdh7rrDGfWIP0YvwZ5DGEhl2Okm4ygfB6WnlN3vutZa/lD
HY7DiEGpoWXCq4JyBwxLAQ2NUp4ZfsZx9H1pAi5MUPGxGa+BphFMCwUu79NJRLdX
UMlbv/9N08tahIev5032d4Do4C83UYguSzMpKsf10mWqL1R6PtfROOr108um1iKO
9wlvtH/1Cz0xSUW04shrkLE/xiSJ9LCw25KF81Rza5x6fcGKgokhK6TgtO5AalWO
2BhbWMHFN2JdPs5GTOpLQ8A+hn3t+UWxg8upRV4JhtJ10TKl7XeJBoqfS9910T0C
ALN+74oKPhbTMU/htrYji+PBdZeMQqu2g1bMva/YspKvOFCrI0Oy6MujuqA5AuG2
/iSMaj7yEvRlZ5ziZaO0gCHIZYopb0Ob9hekb3mhSx/sP8nwoOJTz+dcgjM5Zjg3
9203xfiaweiUJOeFt59zWK/7UYV6Iz3KXB5VeyU+IDYNp0b2XolJOC0dfahrv+67
s7ddbjPSGSPoWdPTWKwrJFW7HYqphpQ2Mr69k0aP05SUgMT7H1aoUFR+rP4apsW7
IhIMZ0wI6ATnF6IimeUGgoM6MJmONZIh7TMS83/GITW0ni4kLkabd50WrMNz5NHc
n+u+MmYQL+xog34BK59ksS3zjO4NjFv4vOtfcJ9RGiPIrnz4nvp7mlfXXNoASvAu
UaC+AtwVAQquSsQ8FMuOf/Pxqyo0Wtn/j/Zq1yxMxWtAAJnHLNMescMrj5oURmb2
NBnPapMgpQ0fLxjrJ2C2kkQnLjwDcrAIZcRUVLiAD4T8X5ziHfD1aghOZ9MVtFvI
7dWRfZwuk93Udu1oySrqc2qKkkBeRKmSFE9XcJvQbzsEuPBXYgoqmOTyAf6mts8j
s4CicgPl2PnrW6J1nfVCCgd5W8AejREEgTr3y3f0hU4FWlopQfmseFqYjj4lK4Gn
4oLjnbrdoI3lcm3F9KAkP5+rCSh/ioaMtY0Hz+brM5kK0yeLwYPe58HuPoxQcpDN
Y4JBnWRjrv6sHEsS8GLT3l4IhY4uJVZ1+5TxITlEfdaGxtTh7hAryHiPcUSWDwq0
vrFueayvZbGG21SHkTsf+drXAGTF7XRi37yfbETK2z2B6yXyrUmqf/821Af+OMbH
AvmJO9D0vXpa8eD1j3YKZLoT+IxNdlatlCPu0qL28onXUN9EkC1Ey8DbqwHBEw41
QLaZJbOpy38xKenCjLUM6S6EqfvnIFJZi3nN3MCMylw3/knnQneuT4mIt4rUrMS2
qYi3UZFA6duRfbr3wFxIwokCm4vMHSVYMy2N0gY2a5zUBpdwm8kSkIN0cQdaSvYA
gmn6E3/oUzvJA6BZgcUQ/1vB77URhLX/t4N/Zsnar9zEoyNpaGMDhUzHB2urckKd
evC75h+s5fz7bpaNbEVIxTP7PhBmPNf+L2BqU1zg/eLOtbJEWXuFi6SELDSWJpxA
2/KO2XjLqM7BlWp8sUoAHRj5FB3iHhN/1Ejcmr42ep3EpJP6u196YTzd17PhD11Z
RXqjAB/QeRfmmZ9Ff4RcyZZ8crmweL7jw8MRPXEyb4JRpis2xP6ScVGaLHP/qiEb
qLo1gk+yZccHF/ftsneE6FWyJUBFz5+E8i4eAkQimN35gl4PbmWvB2JzNZDXdgbW
UMUSpzHToaJxe8FI6joe8nNVi0Il+UV/T5IwSFmveNfMjQmDCN/P0PehoesOJtVq
3OWYe9udXWI3ybu3DTXOU1eIfitoFuTeRMIb1MynfaAKF6rF12lRXVvEJvdBN1j/
fSTZjbDV/LiGf29Swd51dQRtEPMMU2EVCjbqvxRXrZcdi/9ZKu2LtU1ZIKGUlLbk
G43Rrjv8wlb25Y5U9wqUMMGDO0QYTpnjz7MLyMFkiGVYXOfmsimYP6tDyYMZXHsV
HEugpLMGXBjwA+16czheXHLIIvjp8csXxLaBYjpBfzesB9u363eOhQV1Zg/XSxFH
hbgSpbAPWf3esRwQqNvNVnyBuph0BjbgC7U5LNx4vked8A9XElyKgZM9W35DzzF1
IiIUd35hJnBX9V0V1lmuB1wC/pjD8zKNqg8i9No8SsrC7WDjltZiYFOzrWtsNCKn
t4TqjXbI6Y0GdU/bNxm7N32p9E9hIwNwyvm8HN4m2ecdoQpAjxDZ+vMQZfhML3+K
22hyubte61IUbt33aY4QjId7wloefJr7NBal6Abnnux4QCoLNY6O/vBSwOgQ0N/C
nNZCUYKyljpwPcljipoDp+FXM9WjhncxJe2xPfBRr+lOzgjtsYUtvCRDy5yGJMlu
L4usY+Zq5h/8XIyn1sODOUXDQQqRCeNEUBT+nEVqAkx638kEg+kfbixgguo7UeJ8
wjeAfqd79mythZariplnHCF2krrLe45t3lLffq/nzxdTYqRWb6kGklCtcoV9ZUEG
6AzV0Rcts24vSyxV4wsxFaHLsKA9fPDmq5ZonnCGAZXiXkt/V4+0QhjzpijiRWpv
PuCZgvYpq8Nu+RxFk5OLZkwr4oWsOJJ8sC9xRsIjr+G1IohsDZspYuPFQP64iqQG
t5x0cPnPd21CJqTnlJ8iZpUXSbT5wSd85gXiTemBnkZk/uYUdPKUjhEXCPJVnc6x
mxmyAkthwdPm89J2Xmz9Sx03Qi6lnxMgwh+EiMcH1qcST/R9UrEUOHfNMzPoAFbE
/0Ey03iVheIBlbveacpXRXredJmVOH4HwHy+o6yzN92n3SZdeaPx8UkoZ5C+8KX7
UwtladGks7vbMSZFh11HY5+2drwVsM1svTianJXph6X0P7Nddc/5tyeHumZGFRG8
/X/PQVjbask0xzODQIkLEZTzCp+6CLqprfNaxrS+jOmdrf+QeMq7L3cwuOKVFvuk
0ER+LwVu9QjtQ3mMoYTZTlK2oxLVObMmwOvABDTtg7fPgHQTnbXxmCa/LAmcdD/0
2HDTfWBvIzcG6iCml6Ihpk3mb3yy/UUiaaPxLH5E3YOG0SCQsrmxvz9eS21m8dn6
UvzervmHXPWw4pV6WC5RthvXJAT0CsCIQYB4eqOYmS+a/dFrkFnOw9Tl/qdabzgG
RSj5Lt4XSZv/Y0JBwRlJgy7NL/0SfpU9yJiZhvceBhEbUnJpwB5Gev6MQ4hBLEnk
AbU+M/qYsFZxcUy6P1Dk2zwmG4Yolr/pxeUKKlI0bk/vkdpCZVH+8NvkmSfz6wm9
G88lGamCZh7evegR3xRsg+sDXIdIGLPRJlE5i9ag4pOSHKvSFSOIi4qqccKf3PHL
x0XK/LMSwDzcXbWq1+U1h7q/Xg1Uxbvh7vwYHRA9/AIQ4I9fklLn1/gTFI5vgR9U
EA/nqoRllzh9PoCnzlDXBnlcKuEfZWccN6/BRm3aZ9V27JAYoUI//N6JPrAYcxxC
IbtI6zkumuw3yN/nWGAbx/yzxPFcOX9k8TkxVmYAGdugh1jhtuFZc9moQHPNw0+T
jSubDtMvLTqVNil4u4n7lOrMeGhD1Ehix/7hEcyk3csBmHef3C3eCscZbVDV+QGS
73V9znt8gv+ou8uO0dajSD0yhn3McPzSXQbXW3YuySJyfhIpry/KGZJz7T4eoc4s
krYojsQ3MkHSXAMkF8qWsd31i+T8Y4vP3ise/05De69HI8nDgOl1W+ac00JmokRx
o960fZN0HinGjHaoAtFbdT8hx/CMCwMTfpnniDjKasm5gchy6FGpEiUKJJZka+Wn
ZoM/R66xJ7bj50E87SzopWHN2ZB/44noAw1rmQwvb4vBCSPMfh1V8mbUvvKVWVFT
DI3igq0KsCnTqpYb+z7AHd2oQ+Vuz0Ho68H0Z/Ep7KxteMmvr7cC7sL/rQCeZMKV
BKJwvjtqEyUz+8BCfvAEo11Ks97J6InMsPPUBqPzI7WjvU9++O14OYaFdi/jeIFo
WEuIkvhaeVkCpb+3TSWj4l7IYcURGMZTS78bLt9A7QDVTTfVQDh3K771ZNA2hqoM
x7p8N1zTbFnNBQ6TQCSQZLmbEgz+BGo8OIPcGliuYmm3EJgyoCZAXY+bmZ94tevE
MhRgS75FJ1CDV6oJxLYH3x/P2Hg5QfJecuqkqNc26HJXr2Nz/H+h88OcyzsC9fpt
SgDn6hUNeD1M9vK3c3jjxOIaswwvqx1ykhHQVfnL4pXzY55Ew05fIr6vUEmesmtg
mnAW5l/xrjqz7ECj7bm9IqK2RPAohcesZ8JM1zGINqCw8vJz7+KPQ0IqVgDvbfXN
siuNgmjFjl9iBCQGGZJYkxjCYAJLk81NzNGfWu6YD7xuAdqMoRSt458NzFy2+Xg0
9IRACzRSLTv/KZdv37RnioCbxG13fraVYWVnAjciRQLx1cCuBaB5Ncv+63FNMU7d
HMaBpwvdJLw+jOzNeTDyr8oN1V7HtXN3eLi6uBS3y9gAlzb90/bNJXgNqgkepbYM
GSSIs8dBznjkJUEtBr4+1cPJ6NlApyI89ivQfn4zBfrGTIN6C9axGHxzKOQ45iyc
NUmX8FWtqPWwnun6FO9TscqYCrRA6D/bLotlYLnpJfbWzepqGyKfkYzDPzbdqQ4b
LwW0jmCFoiAj8mrnoLidDft3nSZwTiAmVJXmE+DKlsWS+C1FGj9IogbkeVOSC8/N
167jytewNFrKg6mWgxTDwflvascRq1RvzBNGBRmQScHjMeTRZW+J/NScY3MQU9C8
GqlosAG5mn9/xXOXXx7ctjPegC4yFG7FohH9APGnfWPdRjHWkXWSD33VTupQh/Zb
wMcMljo0X1+maUO27fznLhNcXtbGYiOgg47RSaQrn9zZwk8ZgNhnqWN+vV5OI8FR
xeYkFA163FmTkNcbaQ5cjQvP3g8G0XLkG6ukF5X8k43J+CJQUf4nFXCmumwIbufG
pRXqQnJ0AZYmZSXbYEIRRPEdFWVyg0olBJl5nhfH4BvjUbi0/37FQqN6CGpSeejB
CtZPHKnBHR3BlKQQKYl7GDo/ynOli6qGB9ojwS+RI1jAj4uE6FPSdzrJ3Wfmd6rs
24XvgfH2hi84PUV2Jhnx0HFiiRWwrxHyqLwH8jITqFq/oe0NKQEFyteE2o0aut13
QCpiD2aIwwuq5SZUQ5aq2m4JYb13zraBaZr0m2y/cSb0dkwpJ7SXEV983Oa+n2FI
M6OpmnwLGZadbQep9ecmqYpOJ6iqoFeoNyi0zkaNYMmdhLa0RTRtxA0fmff2CtDM
hhudn3M9t5BEIfCxLEiEnWSYXWoLA7mgxaxu1Y3Ba2P4tkUCyLYKEaQm2j6p1+FZ
lZGtfDSFRZsKtQ0HLxarLqTc9WPOCFPg7O7eJzMVguCE4WTngoHlC51PsPNj4VTg
m7az7xFgmI3SAjT58dGgxGoGPaYd5WZDMWxQtrFpChvlpqvx6i064QqCHdjtO/RO
huK89l3TafgPdTfiVoeULbznnDEFdDD2vb/EBtDZPSd/JlyaQktbrSaJj6ZugLVp
9QrOS+jqRxS2nOql3ZPwRUqMv61KKz7L6gjKrn807olUNE2ctAz5ZZYzWYuhhvbl
2ntXwR2U2hDz2x+M+Ne/OhIGW9RWYYp+ODPCy7dbG68IUy+k1RHQk/DNCIuAM4qp
LbTO6i/znDWz6nc/UZDpBU+ypfpOVzW6nrthCqZoKBbbAsMPopcS3OSUiSI8XKJL
WLl3NY1FoYHOfouoRnXTCd41uU442euI4ed0zVTpTVyaNg7EplVo0V7c23h/dtt7
z5dT82VrI/aemzHSPIL1duM7cHVbHdQ51my482Ox/9lgOIAghbDewt6ALkS3XouL
8OqsK8S2DAk9A0kDrV/VnFBSAPk8l5z0xmEIV1WxmX291wEhMrFHBQVujtsBHklm
mLW3javA4PzE93UriajF36OgnHxFPexR6WYh9HwV+Wgtl6ZRJoFz5Q0lY6uBEVJz
LI4azKgbxq4LQdjG9kpA96nvibDEnAsS0uxrM5Uy/t9HYjfIcyk5qzEHUJBPQlef
3sdPUr78kJTXLVDJMrDgLf7vIZIOyaJmeF4V22sJg7dcAVZnd6n7EAynzEJDUS1l
YePp6zG1YWl36guI5b1SC/AIaqJ7Q/6NwOa2oElWnJbonYMQaeF+gkBt/KIOJ9lt
AZnYui0R+SvQ7g6TIBJuo/haShFngY2Fwy/qlqTPMEQtxk0ge4QTl3Franak2Hgi
pLG8ZSo6CQldJYgB7M8eVQBf9hjg5YkEHoj3OEpqHzIVKfp3OAHv65rGLqu3h8ZM
DHbkiM87qpXzT4bcBMes20yfiyohC6e3eo01/rosDg6xzkYR5KNpHhQYLyc1mxdV
HLQsj/J6tXV1Bd/NSAUzDpzAUg+tmOMpURssvC4eFsFyNVXPhUezfddZDHsPHzJh
vlG+VXJervaQT50lxRbp4RL4iz01izofTRicbxQx8LYr0tJ8RbyUeVbAMeurRR6Q
womn+ngfnY34PULD6aEgFtoKhGYx+3peI6fltbxhH7vkcBBFunP5qYGydWFC8LBP
iD+iet2x7j39wv3cn8iQo1Sgsl5y5E5PmkeXdBJKHlGlUkZH4sFzGDp0c2t8n7q8
Kw9PJy4JuGDc40jDThryohNcoqMKspzxPQlbq5QdyFPMl4DNNX6jNPoOWtpr/3cd
0k/K/MqzMgV0JTmqTWTfQLTrafHYg+HBULypk1asCUfp+6BemK03C3iQZr2/0wsP
4GvAYTXLL9lgqGAwzaHE54F48bRTi7rvCRqeTWnSDu6gCoSFCpnKpELVQ0DllglQ
UZi7sjPtRY9vHdAKkUDbKetjP9wtsZpXZ0z6g6ZJYaTW2zEyEZsBHOiYf1zm0K/N
KU9YqS6JU+5f8RV1bUSH/ASx2VCGpsHNWsy6rm88L0hfp239vFjyuTEhGY1Ia3rP
y9vya19wXf6nFBWjQzcPFJjw63y1KrCePItY6CjEg3Ire9DcUtUStu5uIKwS6pkX
zFOWAzTyYrfd4wymHXC29wWE0Uc7gQz3qUtppdxJrjFETkLudY2WjZL1xt4elJ4X
n0LEn+UL8pUc2m5xxvFO4C5JjaU4KgcYwm+KLHDgW8Mkyf3uWBPyymr73dpn1Be/
w5qYkOfAiZbnr/UKWGPLcxYoJnqo8rMUVDSQqiqGE6Uvuftq9frUdJNw4lYb1XvS
aDtCEagTICbkXGX3v48re1FD/GORK/nbDN+26VmgsCNucGFC2bYhjEcLtqwwkVzp
/DoekP3Q+EK0zhsLZVVBAV/riOZTj7RaGtkR1p/UywiGLFO1O+n3Vf/0Xt7Z3t+h
LI3ZO3VrocIWz3oTMkYFJKkAATp8PzTP33w3ZqfPVFZPNpHZRcFfrW6RI6W1Z2nR
CD2Ml63eLNC4fOqib39mzoqdsDYYKi90kXW7ntlKEgI5o2xJKj0/6l7LOy1hGpB2
uEtdLQ7GKUjgK23JUrIASXtkpapkwiBae9wiLBlyuD7t6PeXYi0C4RLPvkw0YKS9
KQb7MmwOnjvcyqqxh9BfuMZ06Bj0btdoWm6dPkCuqCfc6fQ5+amS2EkwjU1ryICW
i4liktoFs2CE/0wmXlQ7P/Y57ZAyp1aCCECPVeZkjRKThCSQF9ysWEkWbPa0bF1d
GEwYyGGQwTXhiDeoNOHwoADmaSHUxhk2U0eQQEjgxbBrzqalPGhYgOxhurv7N8KI
uidlsGjuR4sx7pVjQgAoyAcWl8QaTdXIJeyDgET2iaRGAwOtKwL2tnYnuSpTtw9/
bFAYsy98wjLwuNZhCAW4QwJ6tb5hG7tsM52r+btWYkjNoUb1H7Qd2yoXVVwd3nQE
3cswMJiMDFN5M1/7WoUEhF+8y+jW69S6hri4GWuA4XnIY46EY1kJGX8FQXYnAqhR
B64K36AJRL3YhaBmbxOLz5vM1sxUbalzBTqS6D+r0d1mANaaB54WY2Z4CgGq+5Oe
eusGtqtDfmLx1ZCUy1hmcWCBLANM7eaWgwxln/dr3RYVU8Bzsps59n6h6qEDo6Aa
9HDQImnSiDSFrERB1qEsTAhhqaI+hbkquRd26RpOJifW21jehxSg3PypX9NcHyMv
8RVfbF04lMDz6sT2EsenO2Oz+hcRmPdotp/4bPhgGCo1zN8s5iYn8e5SyWY0E/Bx
tCDN/tPDYUOXUclYP8kiCv+hzRGl9LTZv/Sp/xOSNYoviaDruxJSP3qsTvinjY/7
ZvFkd+kNj6mtEBDYYZ4sE5g2ULBqXYZWi0Y+cD7blPV7lpdWopIIN2Hdd/Ka0Mau
y52hPwvRbJN2LeyG5z1IdMBh/hMkZoodnzOSLQPJX9BSIgSbshb16Hd/i3LVTpFc
DtJYahTEpzdwQ0Jof++XF+W5K4CSYMMmO2A8ix8I2npYFAFddDSZFbgNRhRImXeH
AH6auonbzhK2VhS51wTRqP2ZW/ipMoIEUYaQBc710c7feBbWgd4zMfOMh4W14aEM
uc3gXn6u2oaQW9GqAjHtatMSGw7VfC5hyePwdq3ZHUrcECAD/5GuUiIIPDNRXa3F
jIV7oovepEGeCWvodGk8DjIcuOevR48jEEzm1OT46wZPWGCBjDh9uIxY1KE6y5AS
bh58rP2M0STsHvOurSinVyLUWu4ezsZ1fbBW5XGcNd3xwIK/vCo1Uy4oc6Wi9H/K
0Bj2/yFpRRc3fhg5SmE2lVnJqrL3sNZ3b2rvuNpQ6yQdR8qenZMoZ8O2sQxq86A0
X33ompQiSh2rGQXaJ0MD2UNVyAcNhroryz/qBTdK2vcWIOpA1R5TfCDL9btsp3uw
dnvm9tm/HuzvoHNYVmuNLTQalOvPpKtOhTaAAowWuZJyU4a9HY98y92+uBmRuHty
nWWkkno2hDG7oBxH+VLnJwT+yTbAAT8ZNPDR0z8NhbGyr+7qrrVdtnl4Off4t65Y
0GJWQ2e6FWmjBNYefQWg8QUki1uRqK2JI1lhBdAbiY0mnjzWd/ijvoGCCh4NuhYZ
39YkaVnxFWdoBdjf9VGuYAu4LVOad4rK4Q5xYdKsVtMrkD8YZ8kgJP4yC4frquPQ
KAgubZ9wijq0PP8Sy5T2fNSVbTpdTYGFsn+9A5pXpzPKWZ2PU3cbz8Hc+OYhfs3I
GRFEkSH1swF+V+EgcYUBWeePpJFxlauw3KUOdA3cSmlFBuE5QgBPXTLTaJmSiAze
zt+A3jbywJzWz/1mrynTQ2AWjn/ztvJKVbrhnctaIlLY+rCkdidwNf1pKLsWWzzA
HF7GdfeV8WNWqJNPY6Jf1TJPafkPPVT6i4EfbF+AjvXGSkxpS0caDG83IeX32NEx
HcQKh57vayAkKmAwNMiflURCwu8V313kNGA2bg2+6YS9lKx/kUQqZ3qhHIMS/K1R
KILzOevwTzhuAmdFKmuujksZ3z7yg+GvemNz9ycc7z4NewVabE3X38/yZiYA3IiV
0c6SzSH1fabD5MpIZ6e/fyZ3s8QqHsWC1GM50GMOrmH6fPPhQvrdk3ChJabnFKVP
N201qYmkvgQYcwWrpl7I3Gef3+w2cTjI+TpVwNztzI7QIgF9ESYi09K1TP8R5Bq6
BdC6m80xOi9cENTJpSYvn3INvXSPyyzP1NQsNsa+6Onn+hmhP9FnXD59wBVg/Xse
/8iUGKBDAXiQ/tAH2G1T7kktuctlPQ7u1FMPNQHgvMGfUqommd82bTmYLRKBieow
WMSn0KW4UzS1EIYluEcPAe1+H3HYNaWIfm2SbcydNLggb9WyfvzfaLcjzuM7f8Bl
Qf2xNTrM+2Y98r4ix2C6GfX5E+VY2eChQhHoHFIhLoFsXo1r07xld+y8fiVC0mrh
J05walzOxx4KbI5nGsAOxGCRoRqfuKDXvABWarYJOJYVAm/00GbvwU4nf/uJQxqn
E8/20h9HQ+iiOZ0iLvGmjzTBwgcpB3dZ+JFmaNhkZBsMCXX3L45O8M5NIJIKncBr
WLgPZj7MI+FCPZNLMuiO3ZzC21NXL2hnfy7JJnSwvs5IP/9sQh3C2xwJvNZNGA/y
t4cwmyotSXakBLVs+hTg/9nIZ+ogKbJaRYp+6nFIaV+TG4CxHqRsUtxufQkuWCAK
7C5Q1mEgNXntGH06pm4/sAHR9TLphlbCxu+OjmoTIYPcHcsQTQCqbm9+4U3e+Us6
3jCE2yfltUrxXuoWF6SiXT+eMVkG2SJTs3nhoYdwWmUIH9fQt/pDwQzv8pY2DMIn
Ql4Veux9NDkvovlmAvZsKpeg1Hz888pVvJUGqbl+Vz1+8/b3tO/BTNpoAiprIOY1
y5uTi2/3eT+808y8tFnp2UXDJzZCrzULE//EfqSCep2ySBS+o9YaNL1Mv60d3SUZ
/5UaWHLm4fLVAhSnUidUT95MLhpUAhxF+6cEA56OlaCbJBQ7K6gxKSsC9BQMfr40
SdqOtGC+Ll7SD6M6V9g0vWFNIGaJ4ZjeZalptseaNJaqR9wPwmWuLoCBWXuBB8qb
2lePbesFuWl/EeLo6kxmD9pIUOiv0jnuHwrp7LWCw/7T+iyxCAwUNRq0Aj9K5cMU
YvPuaeS6tsR746XRWfD9ExumWiWZLrU7c3OG/eBTiT+lX4fykMjrFc1oOFeCf+d+
3p98OO0JYcRWbXX5w/kBmquurrf4lc5G/dF09yNnhiPXqiJ+KrYuzPrsbVVQi/o9
hITWLbX/QS1lGuahFaWUvSnhfRn3mVAXP9iMx7S60NuoyCiEblzQLs3Yvk7dplir
PsUGTLbOAJi5/usSYDmNsqEN4mJncdjGpI6A49U6cdBOLEXyN0Lu9HuG+ngdm2Cp
r1B4lNP97VKDjA0VGN4IzBsxJRiEgWCOfHS2W4M6DzN5bUGdoUUXhQ5wFw4M9fti
c+qKxs48FvfIfrYqg2xNMTo6wgbLAuun6qcaD4T54804EJj/HTpzgnyBnM8wezxM
0yxkN1xymwWRA3mZgsn3FwcHbR3U0qWvt8/AmBsb2PYzLEy8wZxZtcwH5ro5G66F
5K29yZos0KsVLhU02gR8Jn/bf0EAT9+PRzirM0nshiiLrXFK7FMS2T3ZYiI1PxEn
0LU05xT3re0ox7l4yqrfEqAgGEBUIc8T0ET9sUeonx+GxcSkOcUlIiJk6n520zNM
wdTspZMJ669JAWStVbCauGFcMI/OoXl6UxdTUSvXLcHk6r1SYZivJiV0WWic+4FM
6GVuSxSJs7Y+Q/napezKkIbiP10SrLxeBO3BHUqGvUdEwE/kpKoDULvbXnbwCHHb
igmqGeG6I0saXfIecJcfMF/QXw/cyeOJsrsLbNanWLVPvxSTCA0o+qPPaMQmVY1O
6mZSESmKdIwYAZ51xQ2LKIA+8T6iIouayy7s2yEgKtU8juBoDQQAf+ZpAgGmi9LX
qHjVTxXrehrm3nzS6xw4tBcZABaCAnkH4e8CuFUkY1DVblhKKD5Nlfkax7u+Ubmq
AHISnWfc6oWIscMIV7xWHauTMr8r8Gs17P7Szag//dnIAOR04C9u2MhfWe6PHvet
0EEhpWCPfwEf0ggzMArSFgYuG2iaxD0leKK/hCLk2hOfd8VvPGAQmZtRQAHJqHOE
p22Es/KwZ5e2cjKxHhm3+CQ9rL2+3l5fBFxbwUABmuGJ3oe/Wzk0lig2TJLYh+yT
ddReASRIBljN1K422tZOJyVwai3iY3UyVJHmEhvIpQ/Sy+PSE5qKcVseKIGKf6vi
FhZcjt4gfiIlk0o408UhpMhX6A+jT+WlIBDGB8H6ws6CdQhtdBsbq+K+GxOLPIws
HIffK7MUOj0Y9haGG5CFGTlyA7Oc8yRv7h/wiPUJb49HqKAptekTNSKHACvGHF8d
FmQAT/aabIF0iYgsuyUsRZNC+H/G9wrSiSz0O+vGC6GSKKQSXzfj2gG5uotwr+il
RcmqjeZerD0mKD6tUZyJZFgoelS2lbmRZKoFuHGKa8xGROUzqDpWLAM2+M+V911U
GoPWq8KZB/VSg+ZvCN4M+AAs6f2HsdDzmHvUx6t3m06s+0cAQwxqP2Bgm0HHD7lf
5Z2F6NLphw480B3D3nh7TpEoInrh1dISxik64S0S6GvQDfLGv2vtnQTjxiIJDNoV
9qHE44vbgTw2t3j1Z41bDiAOHNS0mD6LYLm2hX5d8A/y5aMvTEg4zO35GEMPSR0L
WPHsTqPEkbifmf0Q3JlxVbhYI1nT+i+05elEG2+LmESMB+09YUcAPwSXJL4zaEzG
WVj0NUZ8kWhuFQzHDfr5CdxA3CDqpFYlkC6+y0hKi21KSK8IYFV3dFYvzEFFJ5hF
557dQ89qXYQuLxMlKjlbWB6PfdE02IXgdFJ7r8ixZux4wnwcv651WW8nX2qCVqJK
fYK8XIsiJiBtF25eoUMPzm9Ge7dH+iLaEZUthFo1Dq/qwzL6qEKM/n6O90cBkW9v
qIW9GQSxnf2fIsc5uRPyM9Sg4so2CNCJmcuJyXcLBot/wBPqiqfUNjxuthgUpduM
QMEBTuWvgbYjDD5ha1aL6zqL8qunl3msyAmifjavEif0dMpySnIIuTYtvJzGypVk
QioB0qMHpc+v3mwk8MWOkOAWdvXPFDz6klFsT6yA1bpdhwrn15aeXTro3cWZfqCy
RAqxh2e94BzBh97dE51XwlGy08+XP6Qh1owAdXthWqrSw/qWTFVCB1xJFYT5YZ4W
r+DV2qsU8x4jw0VOfxuQPCKj09tvkKT8yvass0YjFa0hH/XcNWfkeBwto8YJfR5F
3l8q58wmeXuFDc6Vi/ItaA4wS829LBiS3YqOWImGFnlWihLokt13e+8NWqNMogtJ
GmgP2LGVy3sXLam/30IXYkdQfYif9xUgKRNfv1IwL0kto1b4BkTegCpPCS/v1cRx
yXqp0zI7nVYq0QAId98EwTAxZZ6LLtGBR4K2J5vAiRW8q1bQ0MQotJ2SegZwGGQA
ZnxIjnYVUvCDhPd7ddQ06FeJMnC4ddeGkHur7wRYoSRvp8fCUcC25cGbG5iv/wqU
FzL8MW0NQqt4ypuAI0JMxOdVnv0sYZalPjEnSSigUiZicq7g2X9JBzjXKATTuidX
M6QbCefshEHYOUVULffJPTPzJZq3tWvKE3fbIak5IZTqSBzqLlvti6LyMJpq/YpN
ox6FLFABbdhbV/javW+MfL5lSm4UIPpGLNx/pdqTMR8ie5LjDP/bIGkmaod7J1q6
EgmzvANZPDiG1h5NBf7fjOzqMCOo7lcJYcGqCmjOlUojhkG0gprHGMIOZl/jizI+
DJYo82GQGLQG+lhSd5XiXGib8OPzO+1MqvPKci6k3VsUF/ziAqDZ0nRhFpwkHla1
8OiVJnEWXi5Cc0nvp17lSdhOlW2H1n6RyTBQHaW4bwgbv69/Qcc6M3orFV8uEiXp
zicMj0gRVnDzxrcfiyisCnsxGUvRuMYLyszrAt1YTNV8nQ2/Yxhi7LgXo2Z8hUWr
83lGQ8dFoI59VjIxWcx5LoRUTjXk3bEk6h9mcSkO9qUSuMC6IleIXj0npgEqxGtX
tjp2ckD7/sENooOZCrGmJZarYSqOzbqJpUraUbaOZmYa6u5IOpofsdyZPk2Clf3s
KLn4LG48Xq4sJs1/BVbGX0Ms/HyvX8UhgbYATdMkirNSOLpiL5MHVM8XLM5ZwXpy
zogG9dBVV5pDe395E7WQBjdcYDzKJtVoCW13n/pN+gvmcLRRlOIPZbm0+/2ytGGK
2B3n80P4f69ZeRSxzlWbxy5AIghB3qtH+41KHyXDjQEc7bZzOSA/BJMIAGUawonK
4NQSD8fSKcBXTsqoRGa9nUsMuG9PDUr6pHaeSN1Zu67VPkWLwkQJDnTH4PPB0UJb
0q3DiFZFdqPDiiJV43HAR1L/BPBt9t2xtN8FGzQpksNRRbLNn4/y0vqcG4eWcsPO
z/gTTF7obNawrRkwMQbgWSKeA8qpQLLCjFvTfYmcQeNKA6fZoNWgIVYj3yCKpYgr
i6qtdaug4TIq3FvPZnRgjn6s45e2ILog22yYlWj2+zhBmFGhgdwrSmiPOuVsRdrp
nKmtRtjvIazMN2/tQhZ9djE9d5vfcPNL3WEJUt/yasIwqzque6l9drnPURCvZ00F
rzo3DA+d0qI8tcTPmh4wfVEBWdOCWVo4/9PtF4IU34TBoh75E3Zl4imgc4DpPq9G
2ayt5vbNHwYY/JNrrX3thAiGRVseCAY1eAEl1kX90nrYfWnRTqyRnsDkKsEO3kiz
aceZKeTAN48Q0LVBpotw5WpeB/03Z9+bmh4ThPwFB2uQ9Bvw5YZrezna0/Rsgeed
507pQzt9rxpQD7wFREDcww/yTiG4vckbGYwGxqvavsayawGLPxqNwKp9raWWuVuy
g1cYBHxDgsrmy7RDu1YAwDdpwZlB8W7VIBZTSpNAlIoqGfZmlHFv5du9CAY8pyVc
r8noA2sUWSrcWLhB1R62WAoC8IYkzUziyDA5/5vuIX9mvf/5D7s0EfENJnA99d6C
rFbZwqG2kW9HhrNaCVCh3DIas7XO84IEs9LqGRsS8tA5dtK2bGVry6a/56ZPVPHW
1l4NQmst9aEErXTwhCbDLIQcFSzIbmQqs4R6EXbTfGHQLoVLZxQCfe/u1Z0gs+yc
3SxfiT81ZwUNtyOLogG0wqy45KsOiPJh+h3mDwK+UIvOLZaPx3ZiguUPU/dQpGmR
Ld1YkPtSPZU6EwGBsMhUU3Z19Rw5Babt/BWOsZ9r6ByrA1n89O7sLCa9FzE6OSRw
vzNM05Gota2ewUCvUn1T31JDKflBUlJ6njok+TjdQkOoy3DJ5krvtmQlTUsTG2fm
2FcSOpdQQsWU0qUNu9sz/BB9lOpMv3jE+CZj76oY8MkMkLBOT8PpkaF+eos0vwO0
wJDyt5SQPJfz3aCF2fwzxtELu0unsmDaBSCZ9pbciJSh8xGIRWew4gaqnpKaAHqw
cdH2iMP9GFFiqDERAGjvfnXiUXOpK3eu2aYgpMA9xQz1AqtYYQP6H7U0s3sP35rm
CfKWdMzxFe18VsjiUpsrjl0oUy29fkKsXv7vHVQafmDY5IClggCSKbH9NaNuM0zq
mdTKUTE1qB6JYP6JBTp+lepywHQ93WydLYdMaqyUvC/AKT5X8pSc9w8EjApFqWyA
xTxq/JEHUQqgVRoxS90iqBOFD2a5ShVgzrIvWRfLIZlEhKIEEHMjBlXGA1icwzda
durgHL8KNGY846Ko+pdr5TmyYjkH97JLf1I0yUPVpUQg0K55SbLPIAxtyoDe4VC/
8BonUzLeZyBSq7DoxBN/5Wqc7JgWyG9vbuymJRmp88vSQWlFwUPBDExz8ulJeD4t
/uXmaBcQey+8Xck+tomVDx7Ib65O5MaewUHJ1rQsaPkoWAUP7djOMCZvJvIIOExU
HJe3FXLwZptsGdSw50MtlrwANX9FmSJQnvTMIDm7TblcHqV/F/uerExAVuorwNSn
tqNLO1e0BsOKSNAS4YzPJmk2TQZFsKYOaUfM74VKUqhVWvBFUIh4GG1UbvfQ/FFZ
rB7uO4NvfdUZ9x7xhd8Zb1dLliSIO3Fj7w6Aes/7yvMPbL48eGl8uRn551Q0RCCN
+JIOt4WLUUJogxFxDOLj7+U24CpOu97yZm2kGtW1X7Bz1+ZG/JRyCVHGJsz8Botu
BZyde2QKkFtZTTqzPgIMtf2s3SRqvl3blaz9TC5Xwi0w9ABKjeQ0Xun1gOytQv3e
DOMajyv13TVQa3UMQdQXsih23Ck+4lt8q/keIavGo2omCYrTjMAhigUbpRA7/ZIl
8PUER9i26OtmRuLA2ypq06iqvvO5cWzoxvTdoWXiVxGUK0EhgUuI48VTN7ZSmAbo
TjXkSRJDU1tFMaHvN14txb1okbsFFtfvvMxxRMefwH8qTO5LQTgc5FeUONfJ3bQY
HHXuUbOMmYlFBNIRZkK+mPMDkB25tCunyDeHXg2ujikQq1DJJUFddcBhRFtTlPMG
9CJUea1pX+A4HS/RvYfHScpuiJ1YW0RJeIgk25G+O/UPw2mropV0/+sxeWqubWUe
IYbRQCskuhgMYtb8OuZJyinXKM+5AUmbuJ5zWYXxVubRwRuLDPKosK7oPOYoZMRS
8JEPkucXz7XD8YUohnU3c+2F0irjk4lzLQ6CNIwsqGyRWUl9h/kwSKQcN3RBtTl+
0+afirW+92YwQMDVBTZ5IEFjI2ILFas+lmjzIxVRF4LFzE0Ys1PAo9EcG7blmfUH
98fG2tE7nGq38bfLjmx1TajwVOh5erRwD87/8w1VrHkQB4nzSD2AhOXOu0U5wdI8
K/w4KjerW3CYhuStZwvSG9wkRmGeV3al0m+AdDb0aqgwwckezQRW0wBe3Y902fi+
1rSDsuFVai9zhS5K4w5aBJTSx7/HjbxFwocEYz9qChb0ZxYdn3Iz7E04u9AOS9NB
ab3vaoiVlAQn2eaBSojXYAEAGG1JeCmDj3Czm1A06i3kqzpy4QWQZYIWaGJFGPf1
9d38B+BlyUPbz1o7YwL3zYvKIZToE3iD3Hw2vGZLLHVsxt067FcncjYW/W6Mypmr
8vQlyVcMsGQtnzHi53IGvFQApthb+YcNvAgPJ8H+iW8hV9t6TDb/xKkwTbG+Z88n
xCalo+iRW3DCjxCS3FsmovAKzsPbJ1imrYXEz+oRCC6hcbxM6QJHYaBNXixvLn4h
0g4ODKrajvfCtJO3LHf11tbXfJsWwxbnO2IGY9hU/Sm9gpBIpmpBzp/egiXUP8lh
fgzBqZNivWXYZ+s5yc2bV1S12VvvohMIdQ1FTLpDYaXByl/EmO2F1xlSAaHTrTG8
x0j94Gaq0T28mL8Btc2ZBMZtmRkc6m1+WhEENtl4TdIX/KycJSnVMfFDO7f1vOLu
eYyh1sdawFq+qptimGzVVG9KuvSd+xtG7vNqe+xkiOgftJ97SN9bWAxR0IGWeVK/
KSJkNLzXSgzOHFZmQu8g3hVTNCakHMeuliJcEnqqQSEs0plObSmU1adfvULmDpgP
GE+XQgUUuJyNt2QspJUfv9gaoo/NzCpzawZwswL7uhRNlA+bcRMYC/V3qAnJSGUh
a53pWlrrQbW3S/KMwzWKANyyxvUZT4BaUw1k8VeAXvmTBR+zSA/HhFxXq+hov3kj
gNu56bOXMzJ/hR3DRkxnItxZoMsHKSqjsxaiJOYdnmCA3vizDrNbU4maWWUNDYal
lK6S4Ozyo/Aywcsh+nadTMp5WBWrKYQx6mHJGB8nkwg97GBJzuLtgjm68RVveezk
9E6cSIP2PbyQl4pxCk637r5vhDiCIaCb4F32QEYERuMFQ/ccNk+rCGotOJVfYcgp
+PUgD+BocKWAJC3+K9iKbpVdhQkG4ij/T1hRfL9Xr3n0uJZ09qEvDhAdnJoXUCcY
11lDgdxY68GQGBR2wq8r/MAHzLSLdA1jQssfAp9z/Hh76ZnKwKv5Spkd0AVHljn6
M+tXUCqvh1dzwqMOoOtRLDEmszGaK1Puzxd1E54JAio1p+P5aVGUcCcjTL9EAA9b
jJ5neb01TxOsnRT1+Us4r8JjoBhVHG2jIGOfKq0T0O0nvS6AiXWCqeYlvA1qDLRi
X0H2TtjUe461Cq/aVakT2TYpMgyL0u9hvOfijKbRp39vJGc82o3soYJLNWZYOYv9
FWr8CjjrjTdALvRlx7EDwAlZZPFWuJ5DABzPTBf+OKgAfg8xezgMIwU5qxX8pCHR
vmLt8PGYjYkMBJP41OPILXQtPZL4SN9AGfjeatnfz1UbIzlZehm/plZJlOzYZSYF
21xN7SspYcGskNX3yLSu0dcHEk71iN7PgJHWaSAk9spgH9xWk+eXds1YCROyTpj8
4T39EnbEwE8qRQ2GbYliKuFsMKvrOQfyaz3J2QkhrZV9YvvH9zw80TAk9pP9XicO
zZCYwU1eTUDaJpwVmxIG+h//y1vWLKyFwGgMejE6w8sQ76+J/AousLbSJEQPe1pO
85yFmIAyl+nM/uPhP5VEx66Dj+nfINptOFFLvzcYb0dPFjhWXXXQAW8wYcm2QRLR
QjE3qcgy9a2yI9D/0OQe/tWJU76Lk05vUgNbKz0+VJu3YAh8wqvy09EV9aIgYRqX
PWzVqTCdEoalFXZutQGDutqh1GAe7+DDKPARXo/kb2TsRxPoR8hTX04KHe2H8cAN
mYuCIoCDdnGbFi/lPmBe/9cXqX8xRLHxuH3vk1sLrIz3tJGC4ctwz0YLPSOB6Ocw
RgKMQHTcc5k3tTmtFgCzle1KAAjFcIxq3//bKhzAe3iZSBNbbgyPFT+V2nMOU9Tc
XDgAQDALQRcJBHbtULPxu6dq8oUBIUWuh/AbvnvtVT/cwuqB2hnImycyYSvrbQWL
UaFSPQdvh3FaYxPunqOTAWhGwK7rj3Lzn9P4iPv0Vis2v4fFo4hTLpsiHnVru5D7
rguqcZz4NcpnH6Pb+K4sLD5IFpuRhHYL26hFmVU9zeeQuqo2WLb5Y+GWH5AUJ6f7
Lpnl1kyj2aI8LS/GWbggzuYoNh8gxL1BKPD5yulkzrGFI0HQ5XxilfFbIzxzFS5d
t6rOzxsYu1vw1T2uZZtru7tgr/a3yIqciq7AozlOoYDfyKOc88tgQp1OJ+HCBkJ/
EInuPWJs9Xe6YMmc/fQlqoR7wZpe4ER2kJh+yvRlJi550YvHddU5x5h/e8p0bHZg
/Xv5lsnsr45oZ+xlLzAJ/5+cakZdxeyxw2ZwcvOlbO13J+DVR8Hcw1QSDtE5F5/7
2bWE5E1sOZsSdG1TV4tWZb1BfUwXqx2bZYldXKMfel4JmCC6okooVUjXesyF5tbl
UGPxK99JlTp/M5FA3N6eCT3veoJWHzf3rJzIDSAfItRyRIij5ifgaAN6Nh++9PCM
3kBGzJlPDCUFjfhsA7gTFULxtWfO25TMlbGgGeK0uyDLca2mReHxDXj04LX40VtO
NF3QiHRtzN4xKE/q+YpcIrXrLPv2qDZ2V12ijC/cT93CPpR+Nx6lmM9NSN5AEc3p
J9L8I7fYH4yw+55SDkyBWSlIV1rLuBPpY+RzDRSOYpRv/Vyjnt0AxeJkRy7ynN4D
8vUxZhIhp/UYtiPLz+GhpotsR3zaYE1nt1cmchfpuctOhP3zY8bXNI6u5m5IOdFS
axCtTG1N844skCjnYNH5hPeH2nv2/B66NXzJI8FEAq+ReAHDFB6Dc40NoFX29wRb
rrcyFxhq7zuer239xMAOimTEGlT+esRGWCrTEPh7KiUyiPC2sOsnZWYOmOpy724X
RwsLJarskkd8/2oSRJ5T6G+7uCRVfLxVI8lqn8rKcQ/QPrK4t7LsmYaDn03iF2It
h+WC9q5+PyHM+jRGEetNZBmLQanfYhSvVELs7WS1djnfMBgHYxqLC+hzT36jIIJz
8AYUTaU+7lVIYFvdhMcWrXYTyfnU/VtfTb8ZtZDTTDXbmbPBYZAiI3173nFf5UTh
M7VY86H9h3okR0fJ7N0rP65/ofU1WSRsJ4PNwCdk/eLRj9uLUGT4zPIl1N2bFypo
3Kkyc0/MBH38PyPVoBoZvSmKYq5jK5ps7y1aps87NCOhkfk/kJ4/TFQbCkDCuYtK
ploh0RNHNpJFINvBB59IFrLCojUoATYi3hDEeYFShYLwwEwXr4WY4uXbFucVC33j
DzPpV5e0Tc3P9GUZYaV1RzZyZ0vqTlkpNKfHpyxJObYdPgwz0ZOy5qUDzeAkvmuU
tMUINofL5/cGb190GrDnnFRlZjn8KHfz1Gt9igZuee5mcabcdiy0qtsyr3XSBLEI
SrIeOB1HHS1s3IxchghJigPnya1S3LYgf8oNchOfCGkvRGRYZExD6hr5ig1y097C
SCoYP7scExGcgS6Fm3uMQIGBmuHar8D5PE63eL1lWEpeZHGI4Awe67w91nPlJm32
jrkPh23gkYqu2IyJtXDhyFIFhf5QlNae6gcjJcZRripokrnDhoteM2mNxDXLocgc
s6NFYL2BrJx6+jJ+D6HKBww1U7LIZMEQgkrGIRvFfxD73vyQYyWHky/QPImdTk+G
M+tcZCHdiJqS5xMKCbiEGBecdOjWixnw5hnUj8LbKSExh2uHz0QkvMfmizz4j7sa
d4IDeNuDtxbGZTVAIV32FB8pXSDR20BUV8G/Vj9Rgat4DeGdfSOxt6EMgXA02wD6
wx7LrXC4myJhg7N0u1cgSWYioGstQr4W4e5XHxaLhF/hVJmMO9vS0WUmVdhYVlI7
hVSfYNvd1t2Bn8zL+67HxIEoAyzz8mURnMyo3UL2xVVgj+3alXhwZdZuIA2jy1gA
Or2lzF1KrxIFpr52jZ3zNH2fJSUNa6AnfUDsW7YcVeOcVYhSi4nEAMYEXsqYQBG6
yp308DYJbgSvHZCRAH3rcvWx9Ck4xEkjofh+X3Tv8D4PXfgLPdnJSfrrBDHlZbHQ
uEQwsfcqRu5l36uQ4BlMwCbJZunwNwHpEGwkGm5Mn5G/9ILI0RgChEeDlEUY1EAB
MDSmFFSNAcWvWAm/m/33Co1nKFSZZgAW0OuQv2CYxD8bthK+lXY0I34ydrdh1FNz
AMhJzdcCTXOAalLELI0nEkvOzgKaZtJ+hBF7lL9ndGw/9vj0JWoz79hSpqGosht4
HLROxxgME62J08KcZJ3zEGYMiyudtgovPXaysHgenvgSwcDRucdne6xT5pXgLOY2
qylAt/a8x+f8xEj+6h389YDH65FMtUBdxODY+QUUwsJAsRaNatSvETYAvSD9zQpW
CNR/wxKz6/SI7s5WhmF2afhSgIJ+RPYOWhqpr7Fpjfuxw045ox1pq5jjbyvaiqc/
stAqa6kvA49UX2G0UJ1e9RKFkLfGtVKVkd7VLekLoZqS6r/d2HpwNQyZvUAEPtkc
j0OzZQNaCx2TvKAXq2matJX/+nfbm13g4rqEx54MH8XtmQ2mpC3TsJIOt25/7kHl
F3iiQ680zfbOZfPFofCqf0Yc3tECmVaEz+6WOaWIQ9W1EVINP5zHACmod6uw7tm0
A+rRA+kTCD4AZktaSqNl1fEN09p+wkL8pvt2nM2Lw4k+6GwC/iFRp4dRJpwySoLw
3N8mDOKmc+FignmaIhjE3eW8XgeXA+wYIb/7htj9ipzjYJqRmBxRbrDJTffprnVu
VeJ8Sfw9gRQdZ3dQ/4mwT1BRCvBf9mzC/xrsBg0WqhsSu4PXtHn8ESYVPjnzpN8R
l2JDM4S1Wja1bS2UdfMUO/HwLGjUu0J0dx3X32+lF99Q12TfAmTZep2i9trHxaI1
uXljvfCLRrOejaiIVG9pv7NwdLQ2ZDwHEqDluMyyCi0VDMNO1ZurMdyTU4ZBzDQz
/i34WXXIG+34nJ8Uhzmu7KRFzAWoIx+BwYf3n9q8bm3Foxx6Gw7uhsfj4CeMbrAU
p7kNZcauY8BgN9lghIqZxVp32eWH9o/Kk6bEgF5ykHaRz8b2kFeZLce7c/MAHM3s
ieCYArCGOgL//Wz0qp9CILdW8KAy2Oin6JdLPYuplwLjTj6JdU7eqCUv53X4cDWE
HhMayfKDvL3Q6vaep3Q7qbKl0287TknqSX+nPSY3S+5glFyKICXjSKAWDy+N6aYN
2SaKJZpCTp2iCa1muXKhnHOU2p0aSvvPiY6Id6lJutoui7YrXNquabqDxsV2zXNh
f/B/qhpXHlZaykXOKWZutlmHSBsDAltmpgYxkGRhJbFPi5EkfYOyAwx9CcmlHStg
SmUwDQQ+HC2Z3ghEdGaCyWnbQFZel98QndzCbVYvnhZXcvdUEtUe5TCBSzkTLr/m
8FMq07zGDGCtsP6D/vUt8IFjvOKpeUFKjfKXUwzNWMZMiDjHEupdgZu1SaCjwrvO
qE4YyDMDnW/l1mXEJULgkMJMv9ukgA+aZDyOrNLORMMyHZRtGgEjFIEtTJTGVwlV
qrP0uEyCFMVyQvzG1T9lbWp3g6V0utvcNp+FV++H3OCumgfnwCD6iDNrD+d5idHH
A5UKmBNkI3fxqSf88UXktE+e/XeUw8wyhUCmVQ333v3S+sM6vn6pIbYT4JAv9ohk
3MwgL0efGK5AbIwC1UdFzYXKr3J196srxoJHrzbYLb88aljZzD9maWheH8TG1336
ACianHEQfdJ31XyixIdmhrWP75MKwSVZONO8EXUzkqRtA7ZZIGStUCbPyFtqw2BN
ThU/XpM4lv0mybFb4wRkZ+JT7n0jU4wIy7/B1Ce7VkAqq1kY0j1af7swrV6qgXM5
vvCBT7KJeCasspmctFFjzFBrTC4dQU/SM0gLDzAMQTxWqisS4lzdmRqUghl/QH7U
Qf1I9XWXLbPhmXeqIRCYfje+Zq7RGYTo16WRutFFF77U49sPAHP9r1WajFPlmb7/
HaW0OGo/pifCb24Szg8HAIczCVfOXe7R+H6azr9dM4ED0bHIbdPlA8pDXIW2vtmM
JiOD7U1qVVs35h4Ng61mWMYWRS2LXco1dl5twn5QAvg0UpsoY+QRSzYigLSbAXo/
l9jvdtxeLffi1D3x069rOUQ9B0a13LB1k2ECYVJGRf+iNh07+OhMmVqTmKZjbDGx
50mxJwX1r5eZPO+SPTYqGrLPT9KogrDIBEn6/QL5hOhrzH+JUzLuckKCSSBXWhgi
IdSqn3B0jWmLCIk3aUYMMIs174JCMtxFWCFiC1TtDkeSbS/cxKyhuy4cSZVxsh+8
NsZy+Kawf5EfCRE+ga3KGQ2V49JtqEJ62/mv8w9ZZAdGllydwIB0NGPs7i2exSwO
lXn7C4YIP8cwKue04UjcoF67YMH6DMuRK7YO50QV76xM8S7y6OR4efdj1edaiYhJ
1OMq+hV600YliXKDLfwpk0PNaib3sG7/1wq03Z99I7Saymv2XCiJ86IVwrH2Gatp
kFUTT8dER8gxUuLT1743a2+Vyn+ZWZIVOrd+7p/M++XEsDRV7M0tmukXkbUTWa5X
tWtQMkY6hURToifTrMDSB9CpSpXfnwGWA+DuOUsePxsWTA3QpkAdsrkYxMu8ztFx
CH4jfhyoklH7RPXa70qG83FHT5ifJGRJFh/3ac0jWWuTCEVncRx7hxw1x/5/azaU
hsx/o2UIiJ4+4Ws3D/r6oK9LnL63uWbH+4t7R8/pPq4c3HDGz0MbOihKmWFSxMQH
rxB7qsoJ8LDMkUSXI1ejVWoKU+ZqkemrAyYkmZNMp4xUdFRX9xxAYNwfQdHWdDDl
4D47HCTJmTGpRO2ntxsriulOBkNLHBzVv9yZMLk8XO7R6c1r5/sKnOhampFe9pk6
rGnHUvVV/zb8U1yy0n+V8PnHnv06yL8OKUINOxZi5Y8+yAHtkeJjMSwdRaa9df4E
FGXWBlt+WYM8hnN10aysEPpl6Jxg3ON4mHLb5EC2oxKGOGqD0UmsNYbjoThDt/Yu
P6IPYVn/fBtb17X0h4JMIInTg9pfQDg2weZrhQiMfhgKe+Zheg1b+ujuvIHJl4Ea
SH4EUEatJTwLTDrWU+eB03x8/ZDfvXfkZ+QBgpGIlrZOWVhBJgeRm8oZfMOxmQed
C3tVZfs8xld5u7VF3aIS5m2bZi7VvOsvuiShLdgwzd8omkcpTw2AA5JNDthg8em8
7ZHlvWGcdL8PS3YlVtf6XWilfW2TEVCe8AeaXlHHdMaFz3qKpB6aWlB1LJXVt6Di
nZxbkBvLok9AboGTPAAxJIBB6JBlspgH8ErN04XRqy/AR2gvYp/oT7kVr4WtW8n8
f3f8R037XbptMqTZJyzbQLyA7sp+0xiwehHJFo+tJHrXMqK97BL61lCu3BQ/K+bu
GzojWgJkGeMuobF8Cx2+kWx+HvAle3+3EYD2xpXHBWzHORhMNvIRWeJexRqAUUb3
V3oq8DbmsPWEmvWVJr/wjTUyaRzbEBViZI3rAatqw1FUwJek37QdPgxlKd7TENhW
BVhsK62htGKsiaCaEaZSNtOIfU//aYJZysBILu6fjIkRjH4jSqE1bAOb9uCreCAy
sTezYpM8dcDEvBDq7AjHszCt7qM+L4Z6E8XhyA7XY7fRRrFfq4uE32Eh7D7L6Vbl
KYh+SRkqSWw/acyeZqswkikKih+AYlxQf0ioa+7gAG5DHEwY3igGqoVbZtFxS2R8
P1Ae1gdUqqolsQlrIQbMFyC1CaKiOelsnajvKburyw2VGtW36ivh4rGl0zitxjC1
5PoIMNem2/ikOsftJ0YEtb5NnoOMO9GR+WgrOE3WMWMYwttNttoEg8BQKOnbTep3
z9nH/Q2E+MGCPdFW1VWy9nOTRR3ZM2BpY8Tyj5UGAfbJIXYSdvi7XhgZkTNkh+JN
Nu9T8QNrlIIBpzlkgkJr3t59kNjYkMIdUaYKQyMkW5Z6g13k7BFJmMY9ir1wTUmf
RoT6vfSdb2Nz0P706HZVC1u9sMXj+qdxfBim+KSfH4ZYs+6PbtOg+vlDv3zIxiZO
BLR0rV4ROKuzwlsc16FVjUfa05PNNzKD0lwhLfb5mqhHVQewnnskPIkt8tfe3r71
FFpk1taQaXYd6W3wX4y9csa7U8oiKi7mPfLndSFuNzyeSTy1HO424VHV+Q+HRsTu
Rn/1jrQpejcuKwdvaWsqNfT4bkDbwykbR4BadAxk0DQPcIPlNjXqQFdFAPfJTqS9
oGFlaBMnBMe5KQtHcs2iLfs+nAPWv8nFm2BU8sPLOlczrpBbnwM0Je2zA9f3/kCn
Kk9uEtmHnJkix0gvHzgC5c0MRG9KMS+W7wOLqq+3x81IeEM+Y2uaTwm9BIuVcCk1
WE98dLi3NsHMvcARGwolK2Rh73Z/Q8ePwHimzuYgupQe9JL/u50BXuxWkZSolxtd
NqXHGLx05dxMHlxoDV8BvSxQRRV/yEz1NptfGodo8ewHdlobtQbjC49BRFLLiRtx
spurZmAj5LH6NAuhUfOK9PTZFaxhNFzK6LvfLBVFm/dd8KfoGoCnC6at++gaeVWI
KHrwr/RCWdWH1XjLU5Ih5GmfkYGEAUD5EVOWanDgYEOCA0BAKr3oHuf2PZRCabwC
OpgYqEFN/530sQbFwHEfq4dtiL8sQYtcMESwzVLUhML1zcAQphUw+X8dtftgKvuR
cFhWvKdiocDk8ZxgkkL6C8FOSUtmZG7XmFs2Lcij6DWGG/9zT8cj08adgzLDtZQj
Vm65YeP3iKTH+7VX46LzI5idMJ7Zf6xKXtUSAe1AMZMs7NGRuGZTi3dHhJXnVs3t
JBlowhi8wQLd4UkCX5DVpqkY5hZcn5s9hEH54WOz7iX7Mco8fpv4yJUDxEYgwkuL
7C9L9vfo8Brr6UQhLNQbBYyoueCsOGsDbrVX77Sncqufvrc43f4Hjpi/HuR5WtE8
IEWvJZPIydbFE+K7oS48TSQBm0HndHQASfbkWL1TiGrwWC4NIBSzOWWf3qp+WgaB
6Zutua+9WVH4v/Utmoan+oC0wFJaZV+xKNdhAa8RW80ABzebfKm0HNuqn075x6Yx
1L/lG5L/7VXKqr3qcCO3yQd5VXtnFFpViRU50ieUaKd1KqK5aQ0yJaq+CNVeuYVZ
+kNQ0S04HdxvteIfNFQc1i/q2NPUEcKwjnAAwoMbajFVlZQr0+WgB/hcH6HNZQQH
Ac79TNWZBlKFU2OulWDIZUEmicQ1h/QltHU4VTY/jUCF7r+8TdIVega+WIIvEwOr
fw7+xVkNPMjNApCcdnkGePAD9yusDlshw6wAZlx1r2hfl7Zt/eVvs88asKCvZrlo
UlCvGpixVwMWcblyEgadrS32wtmkCNUyJn50DDGorSLHyA4zF0nVM79JyAU9nb2T
IWTz3mf0nO64PrOvcK4QxP1uhSZZePf620YGv81rSQTZ1sQYBgtCAjlmQRAf5I/n
9a4rfAYD9x5txF1rxnFYSccbg3JHs8MR2hzn+OUWKsMsWRwe9rK7e/r3h0SiJZy6
V45qEE80kakrbXAGMqU3fXU/fXexF54vhwIsARKX+Pt5rMtSPwb/nvTVtrG8Rx6s
ngJloTghTV3lyKBS8Gstzs+c4FT4Z8nVie70HQngLabGr928uB12YZyf5MrTz7fU
9+2OQ1sSy9C+rbknpTYnkFd1myNFt6vSvcFIjStj/UxQb0vwif9k8odqaDxhAAmz
n4At8fx1URjTsWVzBrgC41hPxgzcX8l6CPqLbrkS2UlD0mEmcgWiK/VPf15+cDKx
cszyOwNrnlDSRuEQArFQkaX4eF68QgzIPq5MjsTYFxMWMzhxF4xLMXLRJtJHeCP/
6xCU/ImPR7Byb2+MFxEei/khLqw898ygypPtT9DbURjP5lI4GBqITtGht+iHaiwH
snwq2v/77WKpWmC/smvpnscEvo8BSZ6xj+hOWZIHofJLwJHKDce6CHEes+LU3yWx
ZpXLI5kjlxN5qWqfeAgYFNHYScj3IIOtVdXD9ryvVbiR+p/eIeLpfz5lAvnKxXjA
DUZd7TPlvemOf7HKgtBUnInAI43W86Z7wveqkQTgRo2+nl/YxqtyjGhtOBz/KOyj
WfpFzq19xBIp/w/b4SXw/2Mv5bu5sf5bgxQb0CXsn4/MWAv4dx9SNe2GFAAtw4oR
299iWZiHJEmtxJDhMnUmnJzl7pkjrBzSTuexkqWjRt/D/cJusDOTWghTPm2V3X90
OGUmafvBaV9mW2TEt1MlMb1a6x5ky21Nt7fcKuSaAloud6AEUitsxQVicuKGxzu0
Cj3lstqS0NKZDZa2o9EXCxamlatkDhDDLxe68SA0MRmVdjy+PQiQ7KPI3bg5blfr
ksRPAp/iqTTO9wOqqKis14/d7kp+TmgguITv/ouvFC7tuwZbn64T5iYAMKHjQDaU
Caxwj+MSVaItGEujr+twOs52pFHSjDSeGB1s6s3jCMWmtwwsuRqdsILgyZINocGG
TxxBWRH6OHR1CElnlVQ4QjgykDhp7kvdGH981wxAa3me+f5rImUa+Kh9fiBq2KXV
qA3QJbDGhYko9YZCgLrqpJiQgPNzMxnPSKNZPwrJq/77SbDwVFXbN1df4IjEesoT
gmuDtEXuIX61X5yUxslmjWE33cq41SyR3jBOkZy/W7RT53rY1LcMMdn0/VQ6lBQi
zSuz39v9EvRF93A+fFp4tq3tMkXJFJv0hAzK9a2NNEfHYNlHDNx5om6jm8A+VkAj
JfaMLU7tQ0KxxkR1gTQ3XVquoZx652BoMVXizFBP1ZlNwo3dDSILntohF4YY0Xeq
LnZLX7h2Aw0ap8jRq25aZPQvPpg4sr3XGYmXq+xOAAGocxNM/FXT6Y5cGb4eRdWf
UiBQz2oto+GFuUvxsJCDfHpHvuCdJsES6Oua16NHMZoC7kdgOewUHLcwzjPidcuW
JkgU4Z0qDPiS/Ig//bTtI2jd/IRVBnfewXuu+SiiOY1/zG+JpOuM2p31OOqqkwio
doeEjhLNVBpOORX99tKGigXJLrvHPtiQ5aj8PfET/ZVj/HRoo97jsl8ry6ZtL8IF
0z6Ys6omN+dUDH3WIc6u8+9Jm9JdoX6+PXemT1i8XE9I4Q8Apj6A6nC5spf+t5uj
Fn4WUy8qVvJ0zQFSetKxJ7UAS9HORZ6Mvlj5+UkivY8Ds/P1XD2GAvuFFoygDLXR
cGEW5foxpmGVKEIytjNIqQGPvqVOFwmwsBXIUVgDMjjluHltSZDnzDZ/B/tZsd++
4MgvVMBXrtTSUXrQebNtHgq1CA38lj7qwvcpBHs8yFBLJ/l17wgEySgy+z7SO3Pw
cMB7fjxeMuh/ZYHhnAu72BBHZr4hZd4AwAD0lXEsCpfPGcTbmiQ6WvBa/38ImU0Q
jl4f4W2gF8Xub/ZaoAMwa60D1wQBciFQwOaq83Sb8O3iOkn0DYtMLGvZQ6BqW66o
JR4ISVAQTZKw9SKFm6sv/fBmu2huQ/kd+93bCp7wdVxmAbjeFQFiDZ+QT/LhLVlC
KfOcp4V9dA4lajAUl7Xr7hSaR1/WnLSQ7kFGRMyK6n7xwfQjlp8qIkAxQJIIajRk
kq/WV+dWpbF9olLaZUdVqR85WaTgkycegIr7tqyVkCODw7fAXwguAhyXLCbUFHAd
/7lGywuYxCR6NIB/U3CVavQU3m226NXE7RvQZNuNwtuCeJSOkSizyt4wI1JhRapz
ckAQdoXyM6aOiM0hYOhQDZw3oqWzxDGTLA4taw9aa/b+F30kR1GJQhyAgcwykEvV
DGICarKsHLuWQf8Jaun3BhX2sF8mW5Kp6XE+oyhHaAURkwRRx/33jbd2+TqITkOh
XclfVrjxqeUpzEnKienT8YHWia4Rlns3rF3uLO4o7AEeg/ReZHCNi/lKAauAlvaw
0s0Vn1VGH0NvlG02BtoKZzqbORttRQVTeWHQVwKhF6+LWg2bKk2KV3EwVW/ACCWu
8jxuTjkoiwLWn1QEwt8l/l/alq1F1CCjgbyyzCUFLNBYUZuXydhapwahFcVY785b
mHgYB2++niYSiNn18f2t56MUG6VZ0n/FZ26sqVQ4MBkvCU+eLHPsm+TGFkTWTllM
Imtiqo5JcsDq26YyzRUAjoezm4dSBz9+LbLJwzsVuy9zwDVKyPoQdSJQRWlxe7BD
XqIuaAFt9UigqAuACjqIRwP9PujEx0YoiPfa0+gUyqxW5Gocw+3CdaZ8lXTQjAcY
+wV1uVmKDb+gn9J0bE8qpWWDZZq50lQVUi1SwTtNt60sLr9DX6i8xw4OvRJ6QKOY
3aM2i41TSY2JcqnlsPUA0AJuF0kyCq96ffODJjcCGtwCVg35skkOa9f7V8sgKOCG
CwEsFIWDST0PZPZq7SsvHJSxXGMkTBmzrdj07BRpAKamVKZ9+V6FXwe00MemOK8h
jsGqse2iyOePvOb2PJtVcZHtvqUu7iHcQd4YP5FiqB61lPPle7Z+59nKqUbiPvzH
PwaAlsWLOARb+2Ri50z0inJXtC1CIrD0JjK3V5gQgvfvWTCnlt7bgU8C5pbxw9I+
5hFSmQMTjBGwhgIq6So4MJaQ/8I3N/KbuOR6pu89iw5zUbi35mxiDaUZycQoVrk3
0gRtmJiLTZNGIBXodPK+3eYKGjs2vU2IgJ8QSV3lg6C9T3D3lL6QIqI02VTo73Lq
otpljjp5UuEG4P1iieSv5F0wuzgW1huOFLUjE5pPXVbn4xOVjLC8NANf/h8bp900
tDNY2Yf8+xQEw7QPkZL7E6F47khAVsFTtCBq6fOGSdTYMpPy1NzEFRNT2vcq3aO7
uWQG5w2dCtT/LBG6fkz+VQPofpoJt916psPSDv14uX6LxElPtpXqpP6Dzzv2NBL+
nPvuzErNMUiDfK41TXc2bKXgXLUxhWrew9gEL7LtCNr2LRswHfo8ugPZh10dG3iN
SyIkmvjE2x2zr1m8PnRg4pq8K6udWQ9gVBVXihA4dWXSYF/Ko+uilJvmHhHsxPPz
HZNgT/j5CWSbOye23h3xO5/PIzEJpjAUclyqwhdJTkTyjGgeVCQr2f1wDxjt0819
hg6d8DpZgoF3lOnmtdsqSe+FsuSgS+ZKYaEwKj39N70vfvt86yd9m5C/sGWcIGwe
YXDKPL+1BLlkQrdE3rF0MZ4B+SJXkV/fldZUwk9F+H0Jwp7Da0PY03qAC3nu2Pij
dn5FIGwZWuybJKlJj2x5PM1Ts/rqAPvVP/eYWrPWsjMfAel1UjjuduVFFG2DbhmG
i0GNdTRDMnHep4i+HTVBRjEj4sC6l8yCKlKzx3tNyZIs3kEUTAqfegeqIGG05J29
+QZwndfGaL+tUwjm1g015JbM27SJGpUAJMTC4biX5Kl1AlpHZIxP7iu/X6R/Qvuu
+bXBLT1dREO0PvZyKShXtle+ynp8Uub+eH+Nt+VzExsLQXPDlsZd4lBYMbYuyaO5
oC8ywWdmRd55f6hmlgt2xUUrS11qYYr+ROyGPyPVaiqiTzc4qW9NugMlrJip8b55
jghwfTSmArPW1QDInjghzV6S7MZ+aQgyTl2lCVq5aBKhq8/w6j4Nrntvf4/4lWsG
SUvkZm0g/9qBJgcvpzSse+qVjYdgW0LBoZbvvX2odqEONXnGcCk7onJ4tW0TP+f0
TrSbxjYX3uBt88lv8078xzTjzet8GpY/roqCKpbANxJPoo523jEiWzTqLOG3F/mg
FPWYbryyvMIPOdzF5jYfE9e16r5MNfpQhfEgNSyeF+6xrg+PUpvEqhJM2a0kwwse
R0GjudwjN5iQHWW0tCDQFaumJ4+v7C+RFja880cxnPVkZlFu+CrbV56R6IA+Ho5n
hB25msZuweJZgEMDoG/O3bSp/jGY1hv2VPOi2mQk0dNjFd9rp/HgqVJ3bjHIoK4i
34/OBZadgx3pu8MwGtxH4xZneiTzwPi/ISHNpHYq0nCCzBUTuFQ220/8U42fYVDG
nTgpJYYsMLdBFU13CZ0e/x8haFH92i1tL2apMPGrihagE0NhzZI68v0GRQ3XF+6M
Yibw4vqDcEbmTVSMnXF3+FpEOcjlhTESwQz+vbWeNj50/3mx/OvShcm74hdlP5q7
dVow4Q5l7w2dEFuvauLaxNW2muiGd8PQtRfs3S/5Vkr76QpqAFJeBAXkhi46lDr0
9bIg1IL2dPGIv3C37frxPsDJyMzWpzy+hHXgK/bYrMsEPH03B9hBk2PxM/iUsO21
DUQ5orix9QO/K0Cnvo/krsRpDq8+sYkQFJW1hUaecb/5N7ZjnhxdxRW/iC7KezRZ
1kNn7l9Z8ZtE51oFLd9ASoT9bw+JujBEI6qk4jBjpC01hDLMmTnUa3HLXi3GoRDm
NJo/IYZ9rhRsCTOFcv6Gyheohg8MABCBR7ib7HswCs8kEYJU7OfZfOuaWxgWGPYr
4PyhhwYdEIuHCSfAeorL7Nv0A18lIyLZlfGBWGK/L4qz7c0FFm14SUg7vbrkLD6D
6015i16z83KAHbyMT0benj+5Tp7uY7Hbd4VwH5LvdJrpkI2X76jdpP+Wa6/8UHIF
BWSAsTmRxKB3Dyc0B7yL8y0ccFLLiqHuusfCG07ErHYAhU81evo5zrPloHbYFsGS
Bx9bStx1WSRuLcB+KO8uLwLA3uwF9Io6Xfwb0OCEflP44WOLg1oul4fNjqDP4aCl
tf69kCfPkGpF50M7p08M4KBZJ8OmwPAjyBSHM1ZvCvLrw3U+bF63dHwBVli+qBIk
xvp4DQQEoFLIDPH+yrMhExwGzadLATZaBoNLaoph9+dUusD8yldztP6pG5kB5xFw
1UtmAb7uT9BWIxqY9IQdmru8yWXgkQ5WQKAaqnaS64iP9OoB/tdNeiGvHH98G+RZ
5x1Dd0osITn4+cVnHFmSmAm1oersUp7x52B8FzAWRRdc+AwVQVJlv0gWjFbsI3/D
U3XN5sqB2DaUKYGGG6KplJh/n4UBZ/fU0l4i6f7mI1Y00ZrNRFcUAd1p3tI/SSGv
HwYXmoHK4TXt1rDoBBlzxr0KG81w5QGk2nb1ZFxeaD5Zh+TU60Oxo2GzLb5tNjm3
SwhJcppndUqj0CEBVk9pR+JSPqdO+FFkF7vhdx4uGht4peUSyAKdEH/fBeiGMaL9
P8L2mXNxp9q72H0nS2p7qJMZo3H1WEwubCvksW9/01fFUee8Z57Nuba+owVNDhtF
E3tMjzU+/0Y5SUU6qF+/cl7mQA7V4Z1IcuGs+NhejbK2faUIwuW93uEC6yySwBpi
aK7rs+/cf8fI5Yyr8TQIkvhSU5trTesgMNnGKYR81gNDQ9v7a3iGRYSJIBcRkf2K
SVMR+YOBP3rA/pQ+sJbGq4fsGiLWqOQoPvnbNscLSc17FdMj7nZEz6yGsjjalmQB
w8Q0VYlXeEiF5BWexlFlpzpG7KJfGwt1Zfa3cQNF1tW31PWL+wtWevRUWcZm7HN1
JHkffTJ2H1byy9epgO+3kqDycUHvPygWfqiVC+t5yb/NZ4g5ElP1/ctoKCikr6ou
4unmgyLVDKzZ7pKTCp0CjS3vxQlTKITO1KsuoGP4K/FP2uLowcZNoXbclayWIq7B
x5EmdJi/qim79gVApD4b5BIJFj+Vo7rY3pLuRfNoU3fGI7tdoT1P7CMcUgQdpNiA
CTlskilon2W4A+OBZbu6xBPGCEbapy28rqeyUkrSH7rGVugdk8+UG65wI0dchwL8
gtaTT7U0fZDBY1czJLK2NFIWve+pN9eotCHIr88HjPBHYis4RijtVi7oOSXIz6U5
aCpO6D6RVK8DsoPiSh773lef6HwLQScLc2iJK7Hme93svA/A5AVAyIOFKwNdiDxX
0/JbVfUkgGb+KtXykD2sWGLbUqAerqkoItvG8DRrQ23pB7XuCEbQQs+j6E95ryc+
2r2FCj4XRB4AQVpJbZrFf2NgwoqSlDyw6vLY2AgC/RlVSsCNR6UwNLo4R98PUF2W
fyyr11/02CdWiRc0s4CLSiQdhctTfu/a2edQzwIO9g+vYW+nfiqnm8N4vTDdGcGJ
KqZIZ9Jub5Qo5DLMeLaGzCMo4WPnnhshDz0KBh555FyqsNMAm0AbRKtiCF/udIsi
mm84YwdTScYMFeliMp13lpDN43YAMz49xnTvKkbIJKow3jyyq4puTX2QUiDs5hYg
VM2ovYp9n9h3c5A3MwfbpI63a9vAcpOoQ38zbkL2j1rBfMvR1HRb8fvSV9dUidzQ
+73FITiCWQH8laAmjnw4RBcHbM5kCdbYAYh3xL754eeC3srCNaYaVstPNj7pJIdI
ThrpyvIV7hQKZ9PLDeUHtSZSccNdTSKadegXvZL1ceH0rGd/k9jMGM8sMaiVE/d6
DAGSDNgIzff03A5ojj6sTx2ulJQS12gv0DlBmSdRJu/PfoLbpt2+sPGaHBLRcEdp
Q5YXThs17ISSnwWzCjhO0hMyu5nDoGTcB11rRJHVHh9o9nOYcyAUJaZabZWfcSVy
+RrPWR0d4JkqkXnN1C8U5wfU2N26s1b4gVbm0qyeO3bKzISAItEJbZxk8XF5coky
YqYDcEiMSOUm+rUyT6Jxgr34SA8SQ4bEMLPG1nfg6PSeAjq5m1EqXTrILFHp6+vj
v+3zZyxCNTdclVY2I88WAtVn68vkljGXWBDF2h+k5UFjCsZU+oqJLfDR4h2ox9aZ
UcAeO9CiXAIEh3s8faZdYJmnfHbZDoi0O8CJhvFt5l2jaMesSTplsSTjYcna0sfx
d3osugdW6lfP4E/tIYJsXTktJvszaqXJnJqbFOFP9biYg/EGojOxnAw/Q6ywJYx/
0x5lSGjHUcmyoEGF76ERYmfpSDO7y+ZJSrJ33wRkJFKhXxHqjVL3yFQB1+BEPqik
Mi7doFsYv9JkmFKAhL3PdQEK+QC0hh8qSwc3O9WVnDne2D9QdehzcRA4UrQ32nbJ
FhwzTcgZau1Xx4G+hBAfueeYhWE4ICTNpACiS53to0N8v5tSPA3JqA/XfceHTLhb
qymgaalYHMnexYjR9TN2AAW2moJuxDzITAv2SzRbyLPSIXrY8cTownR5ildGqmcd
ZqXTsxD0s84dsmwzADvYffLCrEzhTuEdqYbe3RPbyyS6OfAqbTZ/ZrfbyxfhH3Yk
YydYODLJwpQ/cGbewCjoo6c3rFW1Qja44fZ8MJoMYiAJap9bhuYgKN0r9Mx6kfWk
3OAedOy2qBe+U7GHtrOAblq4iteHaQ3hul80R/I13EDbYXZ18NFfdWCrDbkmHs3v
a2EbI1ECnYUby+O6I0FqeavuDDnSULgRAJAtCMxz69Z56VwW4A5Cp1BMhFWWrIhW
84lRQS7Fmm+GYZOMnfQCKJFAqsZ8ZirHn+J6CUmTD96AVLRHYpBCAGzx8cdjbDLi
2pmKP4Ip6Akoz5xCeRl8/VhIm8hPXmAbaTWmwH0eu2ZGmbhKIj/DzZFTeFsT0VtU
kDYzqHdm/BXnhZnSryFpOY39P4ha5YwaeQ55Bst0M/cuOusmxUVHwGuI/00+j45m
KsszJh3HzW8Ltl+FWGt0jHygU0nbWY9lH/lGQGP3s/BmrnDjLYSCoWES45c4F9E6
jiNUzQWkjA6JRG5n17HSrQ0djxfjmtgtfaWNq8Pw7vL4mfzwP53lrCXprhH8BNcp
NxEwjgIS1qXQuCzCwJWFmjAT14RRMd+lltojfGYO9ZLg6XBmtKFTMJovRlrzXCBI
TW5d23+T4HLjodDyldrkyYQVvfKPn8nFdqz0M9Il/kT6TwrqsbN8NGDar/wuf5e4
IMpNvSKswbJJIlEu3r5ef1TIsLP2qdQ2h1IP3awlDLibtT8RCJj+PmVPHcSzQLXy
WZhO+4MNpRUuVryCGyOAotj7QymZJr/NpT6JsREupV1VWFjFpbaAhc4mfvRZbnkx
cm/hIFm1VDFtoqaaLrm/IInJJsa8zaiN3l/Hb0KDizuKamnq4pzqWm+WNm1cw6vu
0AaRuVT9fk1/ghRbnJJVJNAhcxFFhzVPL0+aY+C9laln+pn8P4G4W57H7W2vh+4c
ehD6QW1Kr94De7kfpMHSPhv+kVRPDa6ss7lU0xmshgjB95ZXY9K2kouQMd9PmEOY
6kM07YXjjSwfdoQiGE7lJg7JwJGBFZbqVPnS7S63DW5hiYroYx9yaVa5gDUshTjU
hsKnEG/K4GJv9c4sWqzK8EoA9Tn3XIag1wzjp3QUoT81d/4FvYj7LO6FBAY+xYRX
2dQItAjIaaJ/QDO9M8uryXei7HZm7Vl6NDKw/M5VxyKZ9wmlIi6bHVLRgRzN2nJ9
1petinxUsRNlVheANqZzA1pYQwbwjKKsTC+litTcfIrZOTAkLHbqHM9F1g7q0ndR
3njJ3EkP7a/8xngh3XX1gIZIEo4pCoISLovHfZmZUoU78d7t17tRXtQ8Kjmq1fHm
4ar5/vLDt0UwymXx24YvMsy5zUU/TBT6TpqQYQatnO4wGbpJx/X0gQE6kpSxYMIP
TJPfDM6mHyhz+8jg7uErLZkvgyZ/DyO/UnJ1/cMKtif8sIK7p9xiVdRk0/sGvRa+
zjhqXJRs3SI/RUmoc/+ovctr0l+oYFnvReYfbWB5cViRJ1YXOxk/OOFTcth2INun
nl+9dWxkNpDV26uRdE/32b1ye29rZeVZNqK43cQusFY2y9QW1H8Yt29qq+lLs5eu
O4m4sYJiALvN5IicU+5VOWvJ4OpG1//AU4P+fY5WReEirOfsITwJZjJoSq18Vm2M
C286h0QyAzmr8O0crqidRO1bmouV+Q3fRb4hvQoTpL4x4zafbt18rjbCP4n1e2p1
EjXTF/Y8tNe+nV7aUpsSGpU67fTZ3XqyHuGiG8cTH3erfv9SYhlksVCY9uZgqQ73
xEhL6l8fdHOumBETpK1dJOSBCB1ca5sOP3cKUaPAw5glOlJLhCT1R2hoo92xYqV2
5RKbBOGbHL+LmBIu99osAHe9mILNBQmmgsYluDm6jLTvk1aoqgiZKhTv9xvJArga
WZqFGoWFWqeci+FEd5vvd9pePx9E5wvJ7pMJZkbmJ5ETUus77ykj7RughoA7Pfev
gnZDYeqcPJSW59y36mL8pB1HWUx/9dBenzaO2E5thVvE/S0esM0x1geZI1ZAKTDi
8hSfCPsOiPJvLRDkeZMeZyJpJDo1jcEmR6dWdwHf+owbMk158+x4nFDSGCKg1lin
tUTbDTxDqm7qwGHCq+W1dV2RCgune/pWJm8q2nM9gTy2BhLztOCaimtsJ8KcwiR+
VyU86uBlcedTP4KYlMPkELmilboq7zL6pOygyJEEQ8nj3HMQkfzyI1DRFZy5C3nf
3r8Onw2E0QP+WeJBhzBJ02PH5bJRt1a1EhKw2APAEjlDD3aDlc5KXWaeRxeTNVF5
hhlYR7aCP76I+xKYpQZj52Uzq7kZ9HFQhOFD5uC55WMByn7lCSA177qy0WVRqUAR
/+1+1+Fo8AEvG1y10dXQ+Di8sfK44YJlHdpSVtk6r+m9eoWNwuD5Mtn/Sz2SeZCw
zKfWJ0oCLNjdTj2iJelY2/dAArSa9wknVH3zEAbGaiQmCrdPTHwg+w/sinyheknO
ZXZiRA8VaY6E80zZGRAbchVmleayjCElKhG3XfJjPe39FzwLuvWW3lJ/YBabHEfF
NRCUmOE3rH5m3xkT0qbHCDXuucf7pKDz2SZsbBavfcTPioIEjeNWDAV/Z3Jr4S+b
KJSBxjZ2xqT1BhHX2FOZOaDEjgtwKCgn/ZjlsKr6B115ieGYvsYtNe8Za2PEd/S2
UM9LsdjQ1fML8kps0yphy18wcCS9sPBm57xSVPHhhJRzD9FgrHgO3x9NxOZxzoiD
Z8Ev2ySkD2MvRoNm+PK90YWHlJTjyjjlT42Pl5jBCgRVwlrZUQzq0bmOT8nnPteG
oTlWQlgVi0t7U3Eqvlte+ttIcL3wlMVjxiuxzedmcIG6L8/Hznst7bujSsfBSd9N
LwKeX5vDk5aE078JffYC4CUXn5AYO/PfdIVf80ISuGb1GAPKdWKKQ4X1ebgeGvUi
qq53bJYW7D2zl0NV/ORRdJ4G7GeoE3Kjd/0L0cPW1HTwrJaVWT+lw9vkYc9pZ3On
rFFAFqjd6qbxs9MoGHxoStVAnb80JFqmDa05wOqGHfiJV8Zgm5onOhdGfkoSbVJz
9UPQv30EAFM2mt3n/bw/aLSpZR5GXIS88en65XLuPLQ8GJPvPokWtSBD37UfWjTW
wDNUTZDZBlCtL09qSa6T+Roj1eFlxP7UAMwkCl17WzgMVZOG0zAPZsXbtzsT9e8s
UIWAz6ANSrTjq3FOyLyI+fL7DM8YBBO7P282vRF8sh7dWpvam9m/sfQcsU8EBllI
1otubzS6S29F+jvFfbsPDYd/6SLipQnEQxWOi/DB4ol7vliNmz1sc6WMX83qA9P+
M5lBoL4wxlYgGK5lsN2pC9toKr89cmxeBYv7+cbKxglzDTDQVqfIB3Q8gM6WYs6w
OIkh2nFHXXcvZV5gj8MM6F/PG4EqnGx+Px7UgeQE6Zyeua0MQR8OrNSLI+3gaYUF
K020pC2lDXRc80Rzz2RqYg+QOfA3GmZ40qPgls4iw3EHumj3sf5VNxSq3x0PzkdR
DF2LnRHZEvmIdggz9ojE4IqSTtMG9pFenKUgjMZoMtu7A2GOeTdjfD0jpHC3q5OF
S2zawvKhekOMOh2J2I3JfQCWvVqTalj4ke4qN1Z2zHuNce2Rrf89rO71Q846IkJ7
j+TAw7y+9W8N//toWb6/azk6POzrM6p+xWD6hhnN9bLNTdR7BErMntNOxdqgJbRj
qK3hKCelP1RSO2gVEpcBDNIpA9Ctn+T+hqghUhffT86PDbvr2MxOFOOlEv4kt+8t
5WUacNfcBPPRQbYyfLJitkoF2ihpyhTXb8WxthWW1rmGAbfmt+1W433WEe7IjMYV
6m496s8nPTJB2ddoHci1sCeVD61Dyus0PIlw0ul6RwDmCgW/Xxj8syE7j20J1RRo
7WEBh8lHAczp7H6ZlxzmHgCemW+Mw3jBbIKl0ILpRH1NSWI3ZEQlfvikVkO5hDxt
0fxzyJrA6DisxX81B4LfVdxLBRPs/DpfeAxvC/vzxEbDMOuCYSMCXolAFwc600P+
zXVdyNUMpusHJk+FpsvYvQxJv0CGjWlbPGArnrM6buXI8YQiydJDkK0f/laedOtS
XpA9qLs4BbDX3K0BACfrxYGltQohvZpWMYD2P2tvqnI4vEMMVgsH0oR9VyMp5oiI
pzdECCZs5ZzL7hgtI3c3gFwMyjq6idjd6LN9UvUIxKf+X21n2ySFE8QLT5kFrgTk
jmo9TG4ZlT6PtV6tt21l9yHXnubpdXLKEwpjMqZStTrs8wgySqlNebB5gRVRbQEZ
Sd/+EF1IDSkI3oV0iEPJfLwjKBZwDKt4kDg0AUvximfWStePFfcz1P7BU4Wj+DcZ
GVp5BauyzX2ATHugaKmrt5TqH8iAZLyiT2mwmUGxICN7mRsFb2lpCxKA6elk4HV+
UhbL93sYg71Loy4iHKx4Ydkdp7rJaI9jKy9FAhrzskw3OLhkVgYVXJjDIPIMYRaL
nav4JHqTCKrMn8ZATv0T3IGBjbSeXv9Z3/6zuBH/333ekCcAE5UhmtO8ocwS/T/j
9f2Ww5QniBxhnyXDM9XD+xZ1U0SSlFgNo+FEPx4e6zx7j9IA5g3G8dMP1o/5x/cT
PUj3UOas8UhB9n4YkbPCKmKWROA2MSq/TQ5+El23jX0WgRznU8ZAA2K302daDB63
tav/Bkn1C0zlZfYND0TC8n8M6OImCJFPnOWW8MVVlTa9OjLFc/OVuYh0igllhXsX
gsCwTDIcrDkArHVNrajz3y2cwiyD/Cgr7737di0wrlZQe7hnweI9Olxvv75hXKRL
J4YGsvxYaB/oJ3BVkvK+LRTyvJTyZsyMDASab17CNsLuZknQ5BT5BAA1y5AwKj4T
l9UdJgYMtNyOSy/18f+RypN+TQkRYih3nWwY9pVv0rs3FYmi2b63awoJ2tXxXY6y
II1ed6Ac9j2iAqNg0G5fqVwyTr+DCxWpafMK+RTF/Bv2kjorATF6Sibnj+H/kp4A
wfBFBxcu7SrLqf6gfi9PiO/DhydCbVcsUxxGKtk1Fpl2z/hpntV2cpkC+TxKKWua
5coSBdLJgQ/M+xszybcUvam8o62/kTMzDGtWlj9rsND2TrgCggfS5TF4X4Uzec89
PS1qFUpuToRTWi5JFwXgjN+NTqLytGb8L8hR5xhqpWvHYVeyJW2r1WKKFvmVSIi8
ehIByLWNzpgE29dyQCa2J0CeiKh3cZBOCqlrwQkc9Lo3nsAdNr1yv/b5Fsb8VJ2/
5txSLrUozOgu591u7Y5R/J8QT1BrIhC9lB/X9h9WdMQdbCq99MAOzkrULl0QaMvt
f3Hb1yKiOx+WstwVkfzi68RUty8j/SXzK6v0AhZF1BZQ+q9GrLmqGy7lzVU6Ygrl
nLrzIGGcJdtBBnrBpWHSbCbcEtocFBw5loGRCos9yZksLjzKfXA8+rMu+eQfbNUJ
qBBi2E35/fhUtAvwEfskxSp7i4jiFLH+0IudAinCvQ0M2/d+psfMjeaHvSYbVuLG
CLRoqUvp4v7qs9OB/eEzyez4N3+bOrQ7z2c5GVX65/xxPj9MvgxMLm2oIx6TbUYr
zNJObwf5GWHYvb03aDRiO5WXDiN8QgVNddJejlz2pBUQrtWpQ14QlQOmM1jyVLbL
29Wc7iTKxMAQNS4rtpxp5speg7ptQeNK4FYAvwO0gwvfhU8IRYh2Pe3hmzZu8kDj
uWb51/Ln85aq16YcWq0MuDbLyOLyjqQ2YpY1eD7OyiouXZzLJ2fJ2IzZ7kIIfCfX
SnbUaOoxd4bs+ceByHv8al4O2O/Tsd3J2PHH4aIzuP1CsyXkYw2Y4YPXRJl8rYoj
gVdkcnrhVrxdpJx2pXdX8fZU3aTm7B1oCq6HRjvrVtV1StWJBBlsK3s/FEZYS/9Y
PC4Lbze162dtxLcGiWMN1UGh+t4Nnra9luo0NLbM2WsZxW6uk/fybviDvMmbMGVg
GiTJAMqYHlzzRNfR0zD+TkpydRFmQt5dEYjTr65TlyK2Eg3OGfNk4j3oZrLZy+F7
fC+iHLRZ8jQ+UT7UfHaSs1+PrLtRRYay8fzV4gk6RJOtJk0frJ6R3scoqLVLTmHv
8uQrz0OEQKAcVIApwD6Qe4CtFyg9KaiUXl+8nc3QnYg2JXjd8r742a7zzalwOFZ7
6GCL2pXZ5vgcboaeQgSgqufiJOv2HhZf+cbv1rN95apHg2MTwB1O/CQ/ZqAJ8r41
KRvja38UTVptTG/tgDhHhSWj9wfCyT7OKclLVVM/qAQAiCN9ZOUfnfn3Lo0gfZ18
oND0T3OUMAEiN/OeM9VN7Eb3RoNHeLyrnEQ4BC6eZ+1xLBM7ORK1wwXw2xtQHJmu
kD/D2wkWxwGqZn1hBShXyESryz4EP/dZa9BvlsBXIPecwyESWSg8LaCu+tZ4kfji
XHw+QvP3Oi60g0B2xSNoZzBXGxa7xeRCEWk68p8Q5MkwsrrheBC5n/XiS8V67zO7
SGaTg2Hj0SURHz58+njahzXZ1d052Zctkdzxg5z6Hx+INeLBl1m1ZmrTK1pD3VZu
tpZrBZEJ6YX7p2uF0FCUu4F3z0jwIZw4tgI7Afw5SnGe5xl9nvoQLtuRrRXV87I3
0CnBk9CM7FyBIjotWAo7TUdv26rgeCxzkZg4Ky596ytPzjMl1d/kkiTa3jtLDBXf
/M+IbDCcOO7j2cThJiQkFq88BiSRN9yAZRmdo5+pSW4Wi76vszCyVd5ne4n2Prnp
FRCVBGPq8UpHOG3Viq6YBVZUY+45cDi9gOz4s+6c1Y3LSLSoCnspOEq7hDGUvuhJ
j7nWYJz/u2VoMw/hFt+dgynSA1Kwn5WrG/sVoT5jtxCVhY0hNQ4TheKyX1GkSEbi
O89aYOfUc9RFN0Az0EQN7jxzjKiuU5KsfHGxp41JECnUalfWYBFneKXINHD90x/G
waiYXlY9kGfrvWqwLPOKiweoTkiMgo3fFoqwxgF2HS4ODA4D2yDmMlg1sn2YIlFm
Qdbjxq1sBKAEFFlK45vabqIw0TT5q7gRr6xapJ9LMLVahldvSE2KXwsNdMSELCOP
FOUwdabBXAk9v8XZXCLfv+v6CxDdxzaE4tyclJG4/Sibh88D8c65Qa8kPpJ+pfW8
C6U6WM5HBmI7xSCQLYfPIh8sQlJoOJLymmp0iSd6OMTAnEhu4GrYLN0MlrUEw+hg
A783SEnmYW7uxqoVxIUxPKCfilyLYGuYH3Hbuwr0SCK2G+Nk/hb7FLwsGSnDdmxS
UwRvR/i3SnieErOqOJ2mqk5oyDnkHX9pKj3kxtgUkLO3g9v36/1AYPLFpsDqImFN
RBc75NNmPoOl+sdpSUmikcZQyvn5AR6Q0yOfurQfpubVa87zE0hVkj6OE2w4OuqD
0b04GfKhe2GOCjQZz178AgLgVwZhdlPFkm3Z9QFNgf22rJMHKxQbr9oxDqWW6Oj8
fkIvk8iU/q2lC0DD/Ea94MUnJt9Jth5Z1wTOIlucSKXm8q/vvh2qCcOJJvigKs8f
Lu6TdY/DbWGeB3Fc2gu/7ZkA7gtVHUBOLM4vuFSKKYVkP0aNfe2NQHVvkSA8PG20
lld/xdoYSuf8ZfFZ7nA4qjQY4EwNyWFRpNkLUKTInYgpbvoBG41M5DUlwiNdXuzt
ixLAOzRspI6uECAzmet6ysCWzXba5qKtXtFcIdmJ/qvySkg0TpJM6cQeza9WcbVp
ItLJ5N5dklId3CtJFDjfrIgBx56kWPeGL8OeAEXizDJR4zlJVr3dwNVbzcOQSLR3
PLfreUAJInoz8H6cP3YdDGGf9QlxdyiWz6uPosUazgG7ShGWuwKxZkLV0c2EFi9H
T/CYX7Qq+gvVEyrkcmEY3ns+sT6YMTvXm7jppHCpqxCo5uA6X5gmkI1+e9RCWWqb
W+eNDbwDBZKU4fdkfXLJWK3lYz+RAp8DuxI2gmWke30eDGBlstaTeMoU/p7d0yRH
jffAvuu1A2Rd5s1Y8jb4oLjHof8ek5Z4Js0cjts0Jbbyx5NM9oiKKfJeUwurrfwk
kL9HxJ+Ck4AIgCjSBnhngb3WEreHEkiUlmm2ssDvsfRfFHFqL4LhyDleu1m0dZSL
yNS+cwZ6YEdBa3Pkqwi9QF3AmP2UpaEU9aqbNoUbticcm97z15a0116JDB0Mrz4s
6IetTTnk98Ss6YM1VveJajp+6Jj57e5dhzSb0YKGVSVXPTD0+z6u1pvpIlZwrfP5
lrPXr6ENS3S/fBWmPJuJ/tbEQNhUr3oGW7epKAax6ydiWnDgdpZeKQsxxoay0OUv
SlNThPyZYdEKO8XLJNQeBkZdfZHIEIF5NTWmM6VlNFux9futVthdverB6YT72qhY
YnHeJsut7aEZOpjOYB3RDEPnsNwmEUp0TzsuGaZt8ixzPRzq+ZnwGjRzxucyY6kZ
vH9qk1ncO8ZZroM8RMbulm6gsv4Bu5coc5+YwnYjFeBx+Im+/LaW8wfouoqwjiD2
8jQvtwciRt3BXslu2936zixDqzHuB2mjKbpeP3W81ofIkOVtRDYt96OlXUByc/s1
GcB0ObhPaR1p18VW8d/ryncRnhxnc3fem+QthMHPqimq3iBlLU/+f1/s4W7twc1y
Yha8FVzI2QH6lyDgPQijeUTN9eqFgL/ECHIw1YIASXzy7+90z+JO7G33lKttJPWO
Ax8doyhk2N5iFF5gPAavjnUeMJBXphllRK/JPcD6IeeqmDwaU9D6m9xe02XhaVYg
3gkEPnX0V47rZszvYLnU75u+Vb8Yly+SwcyfjgVJIDGIatAQPtckjBCLXn5cx8fG
bVDNLywPBEtWcCFvU7YLSEUVxpKGqlRUb/cEbct94NRy5uFLCAzobTZuVQkkJnB7
hLdqz767yp2L5ASkZZiJiJhm80yjn5CvegHViPTdpQ6ZRb7ULuQLhhuL+KWuuPBz
Mw1ixuBX2grbiA7i35RefpcfJhHmgKOo65dNxfR4EeiSuU9D/LYKN04POMgsT/QE
jc+CkbFuYEkL10r1UkHc33wV8FRDMxi4L9ES6HAuLf90eHbjM3aWNmRpnR/rcfSa
WpY8C3AumIniV6v+6oj4qk/MejTyzSeAQ3D+uDsSpt+meBvrMHH/u8tDi1bugeSG
dCkuRAcR5NCSXeG7T6fcC5y12W3vZBjY0kTamg7zn0lQryAKLou0ThIlCNo8dPCJ
wIZniqmwfozhiqphWQZ52UPsknMApEezysTxxehQ68grrbGcta4UJp3JkHBnODiC
ZruTr7jYzoxWs8pWzAqtWWbvi3rfnPmhGyB20QfuLO0DjgL81mK8aVnaoDk5r4KQ
OF4Z2K9ZEW7h49+NnNlei61GsyZss4LOX3KbZuVWJeQw0ZsIxgEoV7zL70sGOvRQ
l8Gym7xQxbfIFUpqcZ3XnrPRK1A2kFtaTOTZIUWmmdcsZVaNzFiZv0pD2C3FbjWO
X/iBl93dDEFkV7HRxuOE3bQPn9S7qIuk3F1QDWFd2w2YzrYKSF5bykEglP3S35Kh
QlQpYVvagAJ03PESvN3IFl8MFCP1jly+7J/147xJgxSk0hqV5uHpgIL+RU1MCT2I
mAhO29iGsfvfEYKR+8y5pvTV2hW9S45i3iqqhqa39YfPtOKvxGh3kcLkCHVeVfWZ
v5FUZ51V7VAblJouH4/aV5OYyu4mBQGCFSh99DaDfFqVzrubjRPM6zMbj1S0MWtp
SaAEbkG9TOpCM00PyZHuE2TCLVW5ejbTRsj+JtERLMEvYbwzMdyWuf4CQKrQ+evS
B1KnjSuL+WRiWPrF7MqM9uQ+8zYqhQnYXDioz42BVtWfVdup67qeMCWP5hs2Ch3J
9D6gg6pNZmy0TCSRaZMPHmuObbLyhpgw1E0rSZefVIF2keycrLjuBzqMcDphh8fz
dOCdfeaUi3OZlKLgzTbapM/9L27oJISeuh0+v3yN+XC80xC003D22SQf+1+Y3q3e
pWe0NFnFPektc7IwzrVUc/oskueLsjMd8+tshr517KTPnkWy3xYx6zNt2z3Ngvj5
E3X1CbFE/PBOsgvsGR9Am8QJxvwV+0qQbU2ts697N4F3Ua4IJnwjLgBBGwl7n0pa
su6g0J83n27oNkOq3QpKB7vCU+e1c0FVR8r7duay1qekxeQK/UmC5W7FB5GGBnqf
bLHy/DmZqTXp7lZk8hZ21dAtwLNs5IeVBeKoXPuYJ79VoxIwtoIGJ4hZQts5lJYh
0nRwH864mOC7Qsb9ULiA9tFHUyhDt8n1/gLwl/6dAbETiw5LSLTGMADMHVu7Yo6H
stPcw4hmY9qIh5Cs8CWO1FCZAckFsubaIxMJ0fOPaZhCypBUZn2XgDj2PUpnh0yo
ltoXKoRwwUrjTpojgqpEdAur5weeKYL4RnnqsKHYNY8ErtPCOfXxEk/HHmTv1FmD
96a5Yk3NjidSPff5erQkFurRbApFKLO8KCrWB59n9Pra35qsQz55w9DeceVcpeeg
ZogIswIgDrYEHqrwZmVk5QWYPs3WWwVCVkt7djWUOXhU5j41H/s10G3oFouN2YZq
2dyoyntGX1TQ+fMmWS598gL7PB2Xel1937jvRZbZS+56unlB85hjAgoUJ1J6deQQ
DpLmj6TbyJ4pFtSUKQmLzWsmjhhpJYeLVxz/QRgtppuoM91T1/YpBh34YRN3ikS2
pHeA0Pjh50tpOdS2zINr5dxsVRvmrVNi1wEc1sWuaFXeqMwwCfItCtrilNcz41qr
IryPIXV83U1VPBtPyXWQ4kjN81XyzJTElYz14VaM/HeVspOKj2aLd2dDU0YqJrU6
dgUz+Qwbagm4iSht9Q5MrHCvTsqnD8ljuy6hi63z7byUT8AyLl6mZ7P98DXch85I
HxfcbEmK93Vam88BK3I+cXXSEWOjQmQM6JxNK0GWAJi7lu5Oq9o0tgjjGQJ84Q9M
fdpq8h37fW1wDu4EANaWbKjogVcUghgo8z8E0EHDWiyijp3RqlM0CIclgkzpgPF+
sEjjxxIq3pjXUFrNA+7XEztE5VB2jD9CcCxVP5RR44f9EzsrkoemrVrvEUZmwOSr
5LXRUg2eQOrpPLdt8yISLdwExRLrPPRCpvyjrQh+AL+BpJ2WHTm5+O49yw0mdKP9
/2J6i+4NXkfUtbdLRCl2v4oitjQF7HMRHcMS9ZuZZa35xoURR3OzHnfw171f2S19
ff7INFqLPi32UMrNf+IhEE7bx2dSZ8i7B9QeVZYIX8z5YbyKgYzB+69T5u1/6OBI
z32+aay2fsWO5IMMwCtZhcla/TYPVwoGTCxHpJV28RyNIUsIk/4DgRYEdAnlp6J0
swZe8/SRwLxfWKE+66mNNfMP5Bgm2IuNbqE/vSiltvWUT+brC5dmLjPC3mqotp8V
WOqJhfxYFHcwRrleiS9zqf0dcb9lbawSPzXLbPj1orkaA3v8CT7vjAQWsFdgHRl6
SaA/zNLS+Ocs/tEifJGpgMu8VaNgJJUQuDJ0ILURk+wDQVLlMv7CsSOyF1IMXBM2
nssdFyHIzzgmYL5NCAGFyjcI4XlalGgMHcetYfZESx0H8yJS1eTBW17rHe0mqAd3
iYOeojIhE9Qb5vcEwWG0KgdmtmCSu6NtUsmdP0P7L5dp9AkWA4RlWPhP6Ecu60r4
Lt58YPhepUC1C1iX2q9ZJpVvzLC/n6QT+ZQl+xQyC7RMBFWbyh5BTh8v+YbFdOQZ
NaxR0wNFbFvVVwh4CGoJ07oWOwcYK8Dl7jP2yEmXoW65v3RMxq5xGx2WSNAdWEzl
XYtn4HfitO4GCyjKjTdzod3JWfxDOlYKj1fP7ZmKjprSSLlCwORxub7sT/DmVQjb
ZxwECsa6uZUrIkw8JHZ3bA8/jIxFfmFOqOH0wdR1Gb4iqkkCe+qUB8vx37jWzM70
xbKzwz8VrhQ5w/5VGs04bNrkovDTqMHrlpthK0Wyvbic0FqU057eli5Xnc49gkKn
TXgDKZ+v4OjGfQXrvAXUwIG/vletW0MXNOrQrSS9KDRfLTvj0dsC/0N4Yncb+WB0
tZ9NCjgjwrQXEm698GqrpB5Uq4TsGwChz+s6IUPCVg0MD8v5MBHhAvAREhk/CRZi
HMRYf+vDtSrVrD+au9ApxnxV52v2GepdRkB/gYBypGcaPnwCSB/cj7dMOH1Vzotz
cb4jGI+fdntNg/pepNAKg+MC22bWvDxVXql5EeVNoJ4mBUWldeiwA1YKFyb3h72v
VoIQUUHelsfTO/y4AgGxliUF2atoRgtms/AvVqy6HH8hE5zetnxLG75xOBps0sU0
HHtHJh0AinJHq/IrT6ogzE6JDXf8DlWamdUZJNO283Ayprk5Tzy645DX8+gObN5o
+T62FAs5i5Szs74+PlVVHFDNoIpRXOQsFqZ1mG8LM2XER/S7h6l5A+HNrPpofiG2
m6OIICX1i4C2dSzyx6tXnM1Ng6sw9j2p+lFgh2GwZVJOIgwM9g4qNAhK/+1IzamD
FIWzS9XrA6RLrv3+ZR8elzU5csVH2QQopgSicfRxRwsd5bnI3WQAARke5MayFfu7
sg1YL3xQMHMv0w1VOBrw/9lDlXIyrb3blVctFhyA5CPn7/HNn0dhDEL+8lAVSHiH
02htkElxZs6ij5e63e+N2bubwXPtQZapwUacepcp9+RkKa6zA6gx0Cpxp8/r85Pp
NoCw13sHehNWKFc8TozTLlkgAXO6tgKOXYYAQvUCJNiEbzZIcq6/eC4N85YBoTXB
+BdhgLYdnyFni1HLyJiyJOGjVMr78k/1sBVw/Dg2/QsI4c8E7+P+Acbw3e6OSN6P
XzsdC7iK9tA0OMN+n5P+RwSVKAw5MPKBffatOUf4P8f2W+dWpKBdDoiVV6Y40QJo
jmJTGYjt1FO+JILhfYdqq7W7zVKhKuA2p36oxyB18O0JiTQklGJiO6sL7BDbtTuH
3VsCV5YlSxCSvguBoab3qlaiqa/bq7z1lNzo+A15QTy3hVHtHFJpxz0RTQNYk3XS
Tei8bGAryUd+1Smq01WDXg/aviZwyjEs3Emq9Mrwo2RxvzPFSOEfBdGFG3oyxbQq
go2Y+3+xV5gTDVNtApitUbGLD7U/esYFEtLOnyek0NWNNMaZI7mmL4tCsH9AFNF+
NXU6Rx79gAEGn4YZ4dHpQrnNSIbvWRU+9HqLFvwwhBAXWhX6Ornu+2e/ltUhJb9i
KOnHYK/ag7VRqWtrLaXNOIqdh9tUkvB9TlJg0Di8Femu12qSoL3eWd7zFZEvlH04
vDlP9fFaOOG1wKOk+I8sDVF8R7CIq54LF0+gamRK5RWaBnTgm0p9EbRHSILkje24
DgxpwZatQqRQvYPCTbjCbZuCZ2mv6MvwcXGz9JcBY/BuRZPXtyKZUdb8/fWeRNkJ
nhYa2G5I8Rsvsdj6oC7TemBaYTIrLEl9XM3bizMMoO5P5ZsbCE5yI6HWUxCU17sY
wK+4E1j9xF/rj2bMgJVZA8ssGDByCw6gwh2vT8LTnkpK/zk6TVX+uCe4Ftd1yN23
X2Q//jTj+yTq1ViEx2piYx1xEgfnMJQWzCApO5jjdDU8jBri1bywMG7xsqTDungi
AYDiZyq77WmRQWHBYN4Iy0aEu3Aeq9FLI1LmeoN2IMV5Rb/cXHlLvqXRp830SxMY
TfmqzUjtRHHn3XyyFEzgzb/fLcYc5iE81jssrNiZ0pByQK/GuF6PEaX/HE77nwT8
YBFAmtWlDvHKh1hPym7CaEZTbN/zxSMKSk/5Fm66OP/yXyD1UHfOsC78PipjlxlM
jWFl9UAq9bIFJCLAdI1r8Cy79zW3QG/cQtnpxNihjKysZT/zIKuzgN/OJtvgUyuZ
Z0YZsDkUkEQCYmFWJAy9zQDwQU7SSd7HBxoileANsdmmyb8/gFPppcTMb/5SXGPJ
kpyGwERMVFVv9O0/W/ufPvaGAh5+r1Vr18ifIDHo0yR5eyT1M9afsV8beyAd4LQs
djj2cTnJeOT43YgX3ItY8ZrSieowMP8id4+OnogUd6rRYvk4kx7bFovt0ODBv5lK
yaH3Pki9tDUeo0yRgF7gmLahlSCi9oKxNt1DNNYIxpgmyU4Y+8G2PDzVZFKHWn2h
ibkNvCT7X8RB34kVlFMG6Uio6y1jIUkUSfm9SiKTEHCi8m4rikttL++D9izL4meZ
3vzWqo0i4PLGDKe37Kj6EG4UsPcHJU9bH9Wn1ymCML3uLawNgpxIvjELVEmdeqpW
py8yQfTZ5vxjKaKvAg7FNBBOKB8yhMWDwKrSF2iEnzdfVPEJtZVw7fSFG8CA9/+m
BKTS//S+ql90uadXEGHpoBBq3TL9s1aFfucWN32Nlo6gffdBAo8sxku8UE7e9VRq
xcwuuDtLOhx/wyfY8xatFWuwwrruhNHsX9uKjX7JU4bryCDAzneQVYJTfxiOyrWS
qGOsxvrA05kQsHm+hp2ZSPPToHL7ZvGr9w1aXx4POqhhu6Grw8ABzFD4gK+xFUOi
sBmhw4E3dA+xrHUJJi9Ce1YFWW0l+Wxf2jFl+84IFh4skZ5NhBHWYZu1TO7dMBy5
NRx2RzaHsgY91VoWCNwITzvtlxJim+N1r5Sfi+qQizTBdmyJiFaxYd4kCVY6r8Bj
K8lcP4ZAG98uRaotjUcADjYQ7an/sMDSJKXcQqLftQbS51mAV72oCqxhGs1xLjnj
pirv9tocoWH39SC1Vt+uvPyYsWMhJ5A/UQo9t4nbEGGkGLBsp8fySAEaAP85F3QZ
ALDdCBAS61zkqPlJ4y6sDS0JcsCELJra0aCW/tm+gyaG1YMyanq11HoRpe3/teRw
Qy7rpGHCyoShuN+OzenOkWi7nWFLfbfRei+U0UZ7Zt33fJ1J8oLXnm4zu8zUUOS8
WScvWeht+j+P5eP5amAY6+iue7X/rMvMmL1az5ZfH623lclRGp94q1/yruuH9D8T
O0TkYs1jb5w3Fa8O1BmaHydLP9xAzWVi4FLrXEbeidnVJEUNmFgyN1Qdaj3uQnsy
QfAgQFmsU0o9oeMys98JrSTambAqfyrDcDTMChaFVvjIXdcis0TEUrzC3CnNigVN
ApbGQzZ+rg1WWMamVa2nGR9sV8j65FUqqD+5PbJ+O2+N0w8xBxsWgWzrF2JU4VyM
CZoDpI/B9+V+mCffhix9nyJGC1h+4l3ZuC5OYil4YSptxW7BXRgDmX0n75VQJFwW
O9rgs5RwsISFEAwOooIKhIjjCfeUGDNsdy/REkw+G82lwSjjjNqSbJ9Qjxy2AUlK
WZbEWO7cbyOAUxdwPZe/n7vfhorecBcAQmHYMgh44TIRuDDZ2zAjmQ3n6QoBq02A
RCzASbJMx2YHqYUJRlMbfq6TOTcXpDRoLi968CR7MFYAsq7axI8cdEITjHSni51b
b0oZYuxcHEf8TtEik9daW+Iit8Hucdfmz6R6QfbBNvQh/gglmuLXwpnxEHiwbUXb
2a6+8s1d1qCZpNVWhF8+RVsmA3KLsKhRnFGsuNKIYvBvmCL737w1Dh9PfL+o6G9I
3MusVgQIkh7nqsc991/Bn7xkJ5IuFGxh3rMXxhY+Nv/VJPNBSWJvs3VZ7PvgF4v2
woZ/dtRssrIJRKKomI5JeBiUJ87mDyMUhIyu4bgB6XMdcAhsJ+Np4sHf6MrLWw0N
v35pfybcWA9uCFQpQxeRogwr0vZzj0mruwztbgHiReXkAQ2TpEg/tNr0naYAcFC0
4WV7kdjvHnANfybNP4uLp71deP3QQ3qd6PQ3ElD0RLj3xGJlgDQHznxMfdkfFBLI
9MKObUHYUhJdDVS5PDgNSFMBy38nKdJrPxZ7zKBWSCgrjZn33vpppUpS1BPZ8yCO
ItR9jtDqdvX7uCC4OzlWLLjO05XOPze2a3uFHvgn1BkH2ddPMO13GN8PB2AY+Ngr
KUKL8RftjyZYB7OkMeyKG1XnZwUAcq08LA8Sear/uvixnFMMxNV+k6jg+NB4v7Kf
6ma4VIuLJu5Q8PShsp6jfRiDl+NHYC/Ym3XV1PwsQRpTR4khJh03/6PG6l1qMLdv
NCXoE5h9KigTya7TkypQN73gBC8bol+TREHOz6cPryT/MQMdMg/NCExLS9UBHIyF
E/ZnyytIkAdvmA2eqq1qez11b+DrZe1Ikg0km/Vfa234RQDfSFlHCoTF9X7APgyC
+8hs3douM5XINGO0n3azhjLHo+tPwyXkgn3m5+97BAJfrQ5mAT89g68JoMl0Szm4
SJTx1ryPAotfBKrCKckGrOuL43G34jdx2jP6nTYnh9L9Slgh51A8j9bUOJ5pute+
fzloZ1Cpw9jfN1Yi+YorejOCFZzYPgZoXZ/Ljk3r0Q8pd4V7EMeA9/6wiZqY9gVs
Demc4k9FLraW4n6rjGakOOat1yjdzCuJaXQCbiHSuAW5luApmfGMgefG7MktjcAb
K92R6SQuEMnXHNhwgrUK/UhCBFRxDZ6HUEapB3A9ByjxAN9U7YUgxtSPPk8Wswv3
VgvmkMTwWnsiEZRdmwbEv7HXBIcd2sTyqhTZV01huoc8Lr7RhQ8mVhijt72wBuI2
Tlcb3JxyzqCGUU5RjpEB9kHaQd909gEOEvGKnt+wog8HOWBjjdhGk/6YfQvvNEit
ORraXzURQ+H729kVs8OQgNZ8MvxCVAyfQgG1AcybIzGBHE5reh4q0KfN8GM2pnPv
qi7ANEg5cmtGlEMcCnaeAWR7JAgjQhm8NTPtPLPFRVrsEaW9K24lSzvKJavIy/ki
LV7wWRiDuHgA0jGyXfAoTpPUPnUptexb94+eQT8pt7fKWSfWMP5g79Wm21RjaG5V
bxuSrJb00Jj1AjljxYyNhzfUTChEthYXJqSX0JNp1NdIdaULL/w4GcQoytFX9pCa
9YeiLj81iuZQW2gaOEaDnnwqzKXL0IULekLRjuER9rGs1eUALNEZ3PA4jxoNvIX5
41nf+03oZmqRhdJOr9vOhLLmthuiGdl3jTXd5ujV9qskMFYpihECqtVsKFvkSTx3
bYTYHolwR0qdHt/TmiT6h4bxEv2nIDp16bamcGT+oF8B3nPfh/Rcf1HuZFNdivys
n/t2eEUun/vy/qDthGE2TueAvnixGBSIHIrgX/8n64TuHTIBDTp0IKYxGX5uzVMs
NqIBD6vD57MghFmfg3gdaJjRTsLvFQGU9dG1floevhJ9mrSAD175wJWTKy/xmXO4
UrtxzFAmOaNZl59Dzuv3F+iZMq4DdJAemTEY/Cp+inhwdePzR2skezdleYErCfQz
V01tv8r1NfOTSqGKcwaRkdh9O8RhXkQnlBQPqcsenW9hU47brLxkZLz3hTFxp1kp
Z0/f+xt9iG0YsTxpIODZaX9RnS5rFMcoo9LrWSUxZ0Dova8G7cvoR4VHYUU3E/D4
FJ/ShYZ+OQ5c8SgQmqx8rBr+m+LDEbaR4PPpreev5n+Z/6DaTjd0m1mn0tdLh+oD
Vg8tdGiJsb8H+5wj6yPn8GIvlyzSzZuG0PO51qKJoHKi8C5Mp5sryWOuMedAt8ax
bMjBSM1xJlDQKSYCefIbjAMGnMLY9ctYYDPQAc8mYmxnfBcOED2p9gcvMIIbQWwP
QiSYTi24xqM6vyC66Y8i36HfrnBZ+qfez8wugS0ERoq5wQx7KQar79KLfbUyt0VP
/vGvuk46XLMsJI9Ts9ti3DklGx6+cBi1nl/iT6ItuYgzcA2Nnu+aqY1hTSV4HWHo
YgcwyZ7KfUFrl403zuhXAmu7Tozgs4hjspqM4zCSr933sNpkUv3uzx5eFGXafHcp
RPvXRN4BfML4Qjae5yr5hcxhE8bHNmjaY1xyUWUzE1vgLOP/lq511Z4ah6S9nfqT
0jCz4ApxARu9sfGPvzcewFOMDXquDn+TtMKolVShBf6Ve0vyzJD+msJHJMNZVSrB
82rxKKDqem61oKpDI2WB+AIJnaKk+EX9bfLh53WhP5n9hYXobU2go/2cLmDZwsYh
FtwdAKJlWcukxoYWtDN9QDl7MCk52y3/IGZqFvon5gyz3InG7tOxxbzLREAVnU5c
jkSrn8h51NRSOwyKcLETzVon1lP5wPAoxw0wcdPHq/jT3b/QY11n3y16YkRVYf7a
/nRnCu2Pxy0vohi57MazZuM+Y/WwCztu8KIUnAxRiZJVxUFzwy/ziGLVlb7lLgmw
af4a4oM5vGI/gBrKR3VMqnWW9USn86AizLn0F1qF2cCYtPXYXm+rnTbiENky2VyZ
4Kuj19VmwFAMWSkB3Slcfz1REMm8Ik7VcLhuKatnlGo97IfmJKMirz2Hi24t0w6i
nSX0yekfTJ/0DcGadBVLWCHdhGRrrH8qvcTSTV2dT+N+xLGMmBWYupJs++JMeZnn
0tKGHrSuXm+G3Fgot0BzoGSYkUPRWs+1+yC9EkkGvu/OUdT17U/bFdMoHGoBTAwz
untruR7/TfdBAfv8OsPCSW7XbwGqa+K8rJ/NGKARJP90+gTtIUxn2VZ6ItnsCqpI
7aIUPgWdPulYJkhAQq5wMssl1OlWsvZhqzuuOc0G91sR2/NwWB1l1EwfORD0AaBs
zxZGbGVuDQg+69UQMhY+ZuSnrIwfWGVar+Sz0OwfL1AB2bwTh8w//uwBhu8zfTjx
dmS/La0O5oa4FoOpQZBiEVJeg6+0F1EReLnuAseJJuCxym8qf1xmJqsLRiRgX1Qm
kd0pPrtsaDl9ObKE2lP8Y1I1ZatZOSJKKdGbufKeBkkbOvRUSnA+eCAdBXllhBtR
gB5YxJ4k+VlhJ+YjrLRX+UbhRANOlIEkWFGoVUneGbrsddm/rpUZYHkJBdEN/v7n
MHs5BKVZ8AorGOqQW6EkA1xUVsYr2ixHPkKamuHMOyLpyFfy+yg9BUGvMwgl9Vks
VDr2UFwzIv7W6rAZKd0PdlEyBg/jcoTpEebsZbd7NeLYB5/eq7rg5a9QTLhqywVf
boLuXUJZVjwK6OZseQ5YeD55GlTbdHvrIkbGEDhanH6IWi35pp+mvF7yvurXGgBU
zU137r/1tQ40axL037YmNTM0+FwcdHgOzMHlMbY1N3aXPuiPt/itBxOcs7H+2w0A
mHiM3/LWzcEbg/4SFAc3hUsR437cAL1n9n3j/yPr8Hl6+NSbXgHNeS0eizGYtT7p
2W3Vz/Id4SuMHm7mY8zn6FsTjSB334DZjT86hh6sIrPinbdU5ymS6cXhitlpZIqh
NKoEAZNEQL0KEcnRQtUUm7ZA+qvuiV2gEAZorxl81pJ4aQT2tmUheg7NuQnaQ5rl
sNr/lPQ0VmiuRcQYlpa9jiZ0xVz9JMxFqOMyBN71N1XD4vu0x0wYmJgH+jIgrViF
pTNAOpkD9fCTuhuMVL7LW5987U9++Dhc2Ux4qpjPbXncoS6iC595rxvMPJnAaF6n
Ud0tqcaA4dA1sYbLK1mPLNLRRbOeIYuiZsAn6T/F/ZlPT5TXp1/xb/RFmQtEObxu
pZtagcMjrSgPXdDOSYg+WFbeOxrDc5UvRsOHyDeEX+lvemMHuahDDWn0wglD+ruZ
q6J7FhQmUHtLmXIZGtqC5OtDpJus4lkm1MSHLowCWYyQS63LJN3ZNEpB5qT6+Uq/
vyW2U4XgjmupnqAHXqiJOpf88joeOHlf2g4oOQFo6du/5ckhnQBZVe+vlMe3YcMS
YTujvFMZ3+0oLPo/Tf/2pu+GPC2TMo1EUW8fs3O9+boRGKeQlovsjD4McpzNVtkO
H8DlVLPEMmR2t68MeBtRz7aUp6LvsAAK0tKHbXpedihr0lgLstHR2MfjcbCYyWxs
XWkbROt7AWsmaNig23z464+hH8XpKfVxXtptFmCgaIzvRIT/7lN8YwXaPaDAygmw
nAjZgcu1PSMyHNErv3XEwDEE7qnmyY+XR4GlgNW2xxa3Qp2pLQnvKip5ZafQN+Am
v13TT3tQfJwHHkIgx//NV50Y1iKsDnVm/3aAwa1Zj+QGLklLO9M3OW1+Wal+wtMw
ZbG9/G614PArnHOcww5uX27MV0+zLjh11q5OgUbrVPlVGf6fdMpBGxOIya2wFBog
YVtzGkbjVX81htVefaN/0agzxMAHzijRkN1xwE+JQcC+7pYfHmG3/b/xofhvVrDx
IT9NQQdqZPaPaeID6EdzaDNkhu54hgHvSa/V/5V44aLQ6EAtmORIWMqGbIXl5opj
EGuE/XESRkStDo6wCvI6Be5eo2DFa4D2P9RZfHAG3cn982s38NlAuWHrnHgZCAI9
J0cjBsb/1dnLD21BRdyFxgraeDLB6ZMUAcZIDcgVAWIHbYZ7xcdM53Fztjc1HlLp
rZcKEvD0bHEKUT1HIZ7CDShakFbRvVmgSTYVQkz1J0ih1XAbDgb4+wfUxchJ+Apu
/cbNfkN5w+Ze518lTUp2X4E5BdTKa4IltS8QUXd4/BlnPOeaX28xOV3WbGwD90Ls
3l0lrQLLT77O7Hn+V3qWT0wQ7dQK/fScM9f8MfcbgOB01BuDRuZ68ZK9h26k2Zbs
DJVepUdHiOaMIx4EYExpg8zjid2Y/JKbTjFeBLJ2GWlzeJ75mdnEgZLlFGnzb6KJ
C2Ue1lcRfYwBuZw20m0nhPhniK3HizRFdeGCWVzac37ypP3g/ZjXVtCp3XjDDbIE
SDcIm3s1FBXB5gXQ13G8JkPsPCFGgz71OmPwcEpKbDyIjPUuEil2yGCvQlilQw+v
9Gz/u3oK7e+yePPZzt2Oi2ZpJDpgNiSMk/drBC5hgTYOngis3aTzBKX5sPzkoPgB
9SpA5HtcOOv96tiqaHh6ko9ULhpGOy5DeTnlg8QBrPMGUfLEBG06vSwUga6dKN7N
/LTFmWb43fyjj+93LBr2b253hjRNSvVoeHfvh/oz8loLhTJXMKkUk5Cr+MtXW01g
hars6Cxkdo/hpyC95v7hfTtlihZEmwDROaZqcy8HzqXhlxNghxWQ8Cmf3ltZaOfz
yfUMsvXK3zvmW+ZS90AycBsT/nXxNLyWn0mfrxJcLXoBdbyFJGOZNTasWqPE9OI4
cNmdK9O2rs52zbJZ3zX+8r4aKu72Z7qFfOeGxpVSMac6Y3SDcIGeiqe6mZliB0CH
xlBloKcXC2UJWfCgOX5cAexb7MPRBtrQnlnQH2qAsClZiCAi2IfvzFZ9TUpfr9Ke
T2ZzdNeg21MUPK/VA/pj9UqDM8JOReb00nwvoa1gqMnA9qYnPyzeSI1RMon8s2Xk
m89I0fyv0lHbhADCKaNrD8xKNYCzQDrcZ/2VcW+vsd6KMVJBaRVxo5/OfjfNbkgQ
L1k6DYbHLFDI++Qkz4mEfIj+yCD3OoayCEDAguS5MwOB57FDMr2D+u3LP0iIajht
fTpGLqTiwuSHYKeFL9YP5ac9EYqNcQtn7kyUZf7lg0GWgshU9PTLv1DDy6gqLVAt
FX1+Zy59tmcTF58KIf25HhHKiHw4NiEimA6QN5XFDTqivyVi/MmUgK8MywDfeaLI
Tn8Kabrau49V9B7QZuT6absyDQc6p0RXAgV8fbD0OXh5DZ8MeionAjXY7yBeI4iH
QAiY8o4U5bP1O6PLki9W70MN861CSfC4HmRGtNyFES96mbPY/Ja6CbeFz51wFJjs
5i8FgY1AqerImy6tOBvH/BmbMDT6ujaH0EjC3HIK+9TdCfSeHE81rlmiEeBzhHJK
C6kzFhN7T49d5y1HlOrxrKwMqoAgNk/z5NkdtiL+jP3v/+oK3xMmSLgO/eJOIrQL
E5QSdXr5xBDHdeSM3RP0ae4F2Rfm6BNqGow/2FHcGgUN7bOWGopHErjLkKtWbF5b
WCqT1THfd82HOvQ57vkOQSZOa488rIkO2eaHpmdF2C4FeSSOFpqubLzIZh0Ra7XP
moQN8TLA1+L73+68o1IMfyJZ5z6OEf4zTy+jXLyZPwqwY6PweHIfoCJvm8N9Wkqr
gnBLw/ZGU9MOHQBbDx3Qhz84ue4GEZAmgDSfTsSIrTDytyDkHt/dnpDBwb6P9Adb
U7ZkiqvHUkSJlJ21skUXsVKoDundsdOuChbuwInyKQxgRLACUDDW0Z+e9syimHi2
hD8biCeC1yr0cSWxG2GkIY108HqGyVpjYKq3x5L0kVCMD6FDuIPoUczWuyqbulNb
Bw131R1/aiI4hAOWslHSL2HioCur6+AaG2fmA9/IRvjgksMFbolBkWoJkykywzZF
vJegghQMxmM5/0u+dYBoLDd8gNIbBRhYtjkWsNFdRCjvNTmqma5iSCUGLIZ+E2FK
Nof1Mh4lOEEG7l5mz4nN8vZLO/Tj2LclasjpnnE41w9W8E6dGDrTLzBpON5juYia
GJFrI1kKUsl1SmNW0n8XSb6xwMOxOu2/ypPwGBNTc9NNC6alvkAsHp2VYwgaBGth
/uisWyZXfsYlbeFdyQhXIbgu6kvA90OB8Yw5TgrShwzZA+lKJ9J6ujjIPuX1oRAB
GDxC/n3xuWCqsxzUIRphOKW+ZcJLv6actpkELcRixOOiFNgGzDd7DjFzPzVpUriT
GqAVeCseHkwkA5ZYWiNY4rL9JRfLDZuRsBNEB015EODGsnT3X9fa5woM3tUGTLb4
fFkE0zIHSrZqMCdlMa2zM7OBAmuCzIr8HO+JXRPjv/NcKSSwpVL3wM3Pcyt7jV26
TXhtKWDuWOyiRcKQuwccX+jxgNrslf+SQ4vrd7k6KAjleVx1xhKYYVEGY11BnF1/
l+E1dWLLK6NTzFWZsYSYzFmdVY8f3K62vnYowZ+dOz8zECvUuW/VzDXAAV1rwpZS
SdvkQwCMg0XD9AeA6LL6mbed1In+/jyMag2kJrzSM60SWn3EaXOAVYm5XiNlkQzC
utUwF5aQ7PI71SQuMgR2o0TQk18mOGfR5ala9t3OQtCaeC+1VDtDdSbhTeUKo57g
7gPvqkCiaMCXChUXh4f5uD/Ch0BFXysG86WI32qy9lIkfuTyzPdEpMH0iVPrrv+Y
3SGN5b4UYApV/6uwLgrnCFJn7DPvrwLHT+vVuhmXwJ3ZNNDKHoWjkoVamffGlHEd
Hc7RWwyQjEeMilWz9T5uYGfuS9K1dtgyfQc4Kq2AcjDN0O4Cp1jyle4cTcLcrxmR
zL2gmupDHweYQ86OHHAYx0jheG++TFdGG2SGUKXwCQABF4pDquH9ioupUMCI5hUb
y5b2GJMQT6q+PHE/xhyA2dBCZQ71fvzZ89batTPxuopqIJGxrf8qa4YMsItNa+V8
Aunyf41ZCXtYjNAG1dKAOZWcMSLiCX9HA0E2NFAXaUbo4n3MvP/Tz8OGk38fUWjZ
YW/IjjDcU4ytDFH02wZtQEGDrypRZH5ypQKZQzxcRjNQ0z/RYwBb5/pifyKir5VT
BRAwFg0R1t7o3qoOrIPv+zMaKBt/PDRiiYKKgtSriuq+mxsSgd2uv1vEQC0utzt2
FI6oTeo2gv7jXcfQvxvkANBMJII4mtGV/llOMpOsl44v3z4qfiW7MjLKYls7WaIe
aBQE0ZblRarb8LMYHYSqgAHBlzh6W61XdhQmu4SZ2bFjVdLJIBZh9UfFp1vbp/QS
dU3GPccMsuQJga8Mzme27g5dAtTIhzH9Jj7IB7gzjkhPi40I88s+VJm7V5iPnUfJ
gzQCZ04mfumqey9mRHTlFMxT+9i4Pfr5Kn/xSxdsc7bG8y+x0v4jtLj2y7AQMKYz
0kTMUKrhI3fk4QlYwaorSFZwJqvW76zPDJ/ZtvEBrVj/muCtLX00Z/Ay9W9onhUe
Um35Ll42i9kNkvoDjRivwRfRm0wrJ+JfNZ8Fxa/wHzLcQJzaOrTMHitC5Uc+kHsp
qz+z1qUv5AafPp3dO9uwxtmmlt3Qtp4JlcaoAEGBOtd7wVUTTB/CmixPFmKXGu5K
3QKfl6Jyux7qO0UUK/JDjFadDDC10kM94zhD3tsYd3zeu9cKKtXnyveKIyNDqWKr
TQdMpFytVwmVRAsVNtcGLkI/aWehVLnidaTqMswI2hWU9fReJX6v6t4VzYv2q/cA
h6rTTKVXKRhd+3YI+OgKbECOjOOILNWD9aT5WZVqUulT8DIbfFkgie18uAxQ6ySd
02foB2vzLJZcnanodkRnw1u4wV1X52IUCr8PvVvOp/KA7CK9xRagC8uaSsHDIsSJ
1ybhoi/jK8AGFoVRMQh9RnoOkCCXwATchzm6Z8eww591uEPdXYMYAiD43ttJ3Udk
5B5kbbhoVUGMupC7KE8eUT7XAuGR44FIqryaPnwi9Vqcx6oT5lCtWBU0/rmigojv
EeI6ldXYskq/pAXfIam5CEUshYw/cgv/F0+ll8HOBPfj2oTRJolA5p0AZ7XeUPs6
dh5EddT+EFrm9pkKEpnS8N3/H99HEXEBaI0hMlTU075dj26T8anX1sKtWhgrTXWz
hUj1v2Ve+3PtY0KKMPU4EmNaO6fStznyiPuaP/zliLiMk3MLhX0/9CHm719TxQyb
A0hImrk2pUQznwDotaGAjzGHMGwF8Px2doBQg1fBpK2DcqOuWOjs1iaYDqLxhXrM
BinQZB+lLDvk9Bs/SDM6htIjzmywXkehZ5IiAqkWKeAtcuG7dS4t8MvFPE3MPKeo
C6Nr1qLVDX9wxhsbKCdmUkw0KelOGqx/hPa27fd09CtaqkAGZSif5vVpH9lo+XUm
rNUKJIGbjvQFq3WxDqqUFa160M+s0gAOktXPcP6pX7xXiGUzuqsGyDGfnhUs80eF
TlTUYxHoOFHL+hNqRwafquR7N0bHpiYaqXuqH/6krHP8lon8zcRJNz2InVcqG3H3
xM+QxpQ10VStlxWCcRfQq25wWS8MaAnQVds6eHNhDIXb9To1nyoA92VNCpBs4p0n
HMfKkhWLyXZS8HVTTi9PDIZrNA//TUN8UZbIZmaTj5xdQ6kb30uRs+mzVTH3MvXl
OF67H2DhyOIHnL33qyx0NferIahAWPZpDsvr0ZHmrmnFI41pambYOA6EnEBdKNGn
jufxlHurOuu72CcQZJ4ocyXSYgxk+Ve2tXRQhWd+vGUNGEy9miPKItU+VKFlzLPK
41O0U8bM2GUnbdwXBbvaL51hIiJwdTWF5c8SDZmwCLPRRDIytp04E648q8ZdqK9D
LvsN/tH+ck1F5GF7BxKqV265u94IJwItnEbxGrOOkPLm9UCx74TzSPpYQwpAgxfD
jAJVuFVIuJsv5MMl+fKRqM1lqYVrOTIbncHuoZcWtjgt5co3bPvPvpS6tKT+VMj/
HuiuEZSzg+UTqZPEPWCIcWd5UOxHv1Vo+E+3CehIPyJNNrBK/TkXszygy0W8oGIA
N8HXKR7tuPI5zI9BqTwX6ZvhFeuD5ZPjBKABnTQc7nNQLIti9BuO5L1f2JNZdfrO
gm0z2lMkoqxedeeA4Fcdctpuqtt5C8tTPNtqFYZ0nx0Gz8KuDICKjdaWiJ2r419p
FEHZzlIWlFcdk2cbuCys8wcCPDhuPTIFSYm3bAh422QNhcKtxf6f9YvaBVhkE/J1
qU1SBHCPZNLDy9FYEYUkH2dF1Cn9EqwXVtabd5U4xvK9AuY5doFZ2hDoiXQgavaH
faGuevJGUoj1w9j1I+neQnVEwjfkfnzjVxR1f3ed6I6FvZALE+m+HSCtKJ/ujIP6
GTfdTjLwex0ouEmc2woMlQQhU+vzl2YnYSy1DlK4IWODNcMZocoKIkhCQSdn3Mk9
ng5qOSkKJVkBtP7KEGOSgSHCbdNhXUUeeqW5xE8LTFIl+R5osak9A7RB8tBEq8Gq
uD79ar5WZl7tlEeQgueUkKx12pWsgTFaU3s5Npwyd0bjm09AH/dvPM959Xp35hLL
ST8I5x1rBkNJROVVALm8ZcRl5Xhe13gigfR+oXuN8BXEKUb7FU4E+mbAbUjpaI76
mu12k7aojN6n0CCBh2FA00g/Tf80Ipgh4m1ZwjNV5qIk8kHTvTLdvswYJRGWJEkU
XsxCnC0F3mhgXdYCOBdqdoNut8B1UCZHGmsvJuG3mg3xSOz4wkG4rCuODvtgqjDV
aWUdSPmW/0+PFCsAUL/8bevPVdKgIwuAe2xr2RpRgvGGlMRCXLV/KQ3B8wp2DUjm
936T19oveYVXRFtHiu1Adz9bcBYDWdXz+LIyL9Fe+iBglQD4ao5EQ1DdtlO5oN/+
Id/Yr9tjnNE22td/o744aoDkAO8WXUDWyvbi9wIly8O/FrB8MCNfQT2PyjOxIPXK
vVBTRRou6j85lDDXdrq7KIrY4RqXKBu0V+TkqsxFpQKEi1AgJbEsiCN98PDuq1n2
Oo3OZpOHlTb86UUlICxHWUpjMng5bi2h16+/l8PORg/mZHmAOMt6KeOz0NwPuD8W
QWjFL+RqTp+6+qgFO5sZQXZj+0PZiN5zEufqOHQpX76z0bFr5Kxo5MQvG8zukJZD
Prc6u3aWZf6o+czXleogHCY3UUK/e+0eyjp3OubyOE1XYD4IB60proVj1IuVzKgx
Q8E1XO34QniQxWAmShbMo2dkzpTUOLhHJMZ9CsUK+AXDxlg6fppneyMW2Nw4Kjol
oBZOJbfBlJrCJEcK0PoOqmJOlFSgbX3S9Xgd1XyxN6WcjvD6FarWtfs+wU2vi8Ro
/YIZ72EJm6H9sQZBqFK7WwGbTLN8yadd8hj0pNjn0JY0agIwZ1aIMqk3lmchCqNj
4hrIc8C5bsJ2KMeTnZM8FdvivlbYKVTik0JJECbz31MWKAPiai6uPR768SES//sZ
s5OjUQKA69pxLqy7czg2yKygBHTUMcqICpyPi5LMrt7R16i/wmnLy6s3kkO5TGO6
TqbxRMoTDinRB+J1c+oo4YZfQlXyTcLqeVn7D3LokVa3TSR4e0k8D/60es+pzuBP
hAE9YNBGy2pxF1y5SY+IxeCI4xlHeXiPmhGAsKdxiccrtogdof7zHPT2Tkl14T1I
mHweIViDrVl2Hpr0WCp0uIl76LNkbUN8fT7C2bjRoz/I4MqfpiiiIDPMf2eQnjEW
d2orpDxYOZ/KeIHm2TGE+jsopnFy70UgW2y9TOpUZnzj0ciJv6m/Jyxbac0nh7MX
0iw6Fb/0f+XGzG2oPTFE2QmG+meVMSaIp4zxQTEsMhFiS2+rHct/p0NeYNq5/H1z
eUc5JHZIPCMdyG2Y5JMDL+eV6hNE3VVagU11IRZ03LUhv8knpRQ7DkT8p+xeBpE1
J7eN+6yShgDqSXVWuwrFa4rthnKM0zTYoWBf56K8KW0JUZ8MTj8tIUiyQjmmB1Qc
KJd6t8UhEy7KzN4jxo0l5vAgK6GcoXCn+eh0/MJxSHP0q0ozCbu9q5LQ1dX0XU38
Q8c//I9CC8AJTtFbijMLwLFySK7/DniMI1hzgRA/Ftk=
`pragma protect end_protected

//pragma protect end
